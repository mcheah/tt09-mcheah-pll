magic
tech sky130A
magscale 1 2
timestamp 1731255094
<< locali >>
rect 8717 2774 8779 2799
rect 9180 2799 9215 2802
rect 8813 2774 8984 2799
rect 8717 2765 8984 2774
rect 9134 2765 9260 2799
rect 9180 2739 9215 2765
<< viali >>
rect 11879 36418 13348 36452
rect 10882 2848 10916 2882
rect 12630 2848 12664 2882
rect 14470 2848 14504 2882
rect 16218 2848 16252 2882
rect 8779 2774 8813 2808
rect 9486 2765 9520 2799
rect 10974 2765 11008 2799
rect 11234 2765 11268 2799
rect 12814 2765 12848 2799
rect 13074 2765 13108 2799
rect 14562 2765 14596 2799
rect 14822 2765 14856 2799
rect 10587 2629 10621 2663
rect 12335 2629 12369 2663
rect 14175 2629 14209 2663
rect 15923 2629 15957 2663
<< metal1 >>
rect 200 40607 24146 40629
rect 200 40051 222 40607
rect 578 40549 24146 40607
rect 578 40205 17326 40549
rect 17646 40535 24146 40549
rect 17646 40205 22672 40535
rect 578 40191 22672 40205
rect 22992 40191 24146 40535
rect 578 40051 24146 40191
rect 200 40029 24146 40051
rect 800 39559 24146 39581
rect 800 39002 822 39559
rect 1178 39405 24146 39559
rect 1178 39061 17326 39405
rect 17646 39390 24146 39405
rect 17646 39061 22672 39390
rect 1178 39046 22672 39061
rect 22992 39046 24146 39390
rect 1178 39002 24146 39046
rect 800 38981 24146 39002
rect 800 38980 1200 38981
rect 13637 36816 14062 36820
rect 13637 36764 14000 36816
rect 14052 36764 14062 36816
rect 13637 36760 14062 36764
rect 11753 36572 13361 36592
rect 13489 36572 13606 36592
rect 11753 36452 13606 36572
rect 11753 36418 11879 36452
rect 13348 36418 13606 36452
rect 11753 36412 13606 36418
rect 11753 36392 13364 36412
rect 13492 36392 13606 36412
rect 13635 36218 14060 36221
rect 13635 36166 14000 36218
rect 14052 36166 14062 36218
rect 13635 36161 14060 36166
rect 2031 35093 3068 35099
rect 2031 34987 2047 35093
rect 2535 34987 3068 35093
rect 2031 34981 3068 34987
rect 200 4181 16189 4197
rect 200 4175 5058 4181
rect 200 3619 222 4175
rect 578 3619 5058 4175
rect 200 3613 5058 3619
rect 5122 3945 16189 4181
rect 5122 3613 5786 3945
rect 200 3597 5786 3613
rect 8829 3136 16189 3945
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 10870 2882 10928 2888
rect 8763 2862 8883 2878
rect 2031 2794 3494 2810
rect 2031 2788 3330 2794
rect 2031 2674 2053 2788
rect 2616 2674 3330 2788
rect 2031 2668 3330 2674
rect 3478 2668 3494 2794
rect 5039 2751 5049 2803
rect 5101 2751 5111 2803
rect 8763 2774 8779 2862
rect 8867 2774 8883 2862
rect 10870 2848 10882 2882
rect 10916 2848 10928 2882
rect 10870 2842 10928 2848
rect 12618 2882 12676 2888
rect 12618 2848 12630 2882
rect 12664 2848 12676 2882
rect 12618 2842 12676 2848
rect 14458 2882 14516 2888
rect 14458 2848 14470 2882
rect 14504 2848 14516 2882
rect 14458 2842 14516 2848
rect 16206 2882 16264 2888
rect 16206 2848 16218 2882
rect 16252 2848 16264 2882
rect 16206 2842 16264 2848
rect 8763 2758 8883 2774
rect 9474 2799 9532 2805
rect 10882 2799 10916 2842
rect 9474 2765 9486 2799
rect 9520 2765 10916 2799
rect 10962 2799 11020 2805
rect 10962 2765 10974 2799
rect 11008 2765 11020 2799
rect 9474 2759 9532 2765
rect 10962 2759 11020 2765
rect 11222 2799 11280 2805
rect 12630 2799 12664 2842
rect 11222 2765 11234 2799
rect 11268 2765 12664 2799
rect 12802 2799 12860 2805
rect 12802 2765 12814 2799
rect 12848 2765 12860 2799
rect 11222 2759 11280 2765
rect 12802 2759 12860 2765
rect 13062 2799 13120 2805
rect 14470 2799 14504 2842
rect 13062 2765 13074 2799
rect 13108 2765 14504 2799
rect 14550 2799 14608 2805
rect 14550 2765 14562 2799
rect 14596 2765 14608 2799
rect 13062 2759 13120 2765
rect 14550 2759 14608 2765
rect 14810 2799 14868 2805
rect 16218 2799 16252 2842
rect 14810 2765 14822 2799
rect 14856 2765 16252 2799
rect 14810 2759 14868 2765
rect 2031 2652 3494 2668
rect 10575 2663 10633 2669
rect 10974 2663 11008 2759
rect 10575 2629 10587 2663
rect 10621 2629 11008 2663
rect 12323 2663 12381 2669
rect 12814 2663 12848 2759
rect 12323 2629 12335 2663
rect 12369 2629 12848 2663
rect 14163 2663 14221 2669
rect 14562 2663 14596 2759
rect 14163 2629 14175 2663
rect 14209 2629 14596 2663
rect 15911 2663 15969 2669
rect 20749 2663 20759 2672
rect 15911 2629 15923 2663
rect 15957 2629 20759 2663
rect 10575 2623 10633 2629
rect 12323 2623 12381 2629
rect 14163 2623 14221 2629
rect 15911 2623 15969 2629
rect 20749 2620 20759 2629
rect 20825 2620 20835 2672
rect 800 2576 16189 2592
rect 800 2570 5058 2576
rect 800 2014 822 2570
rect 1178 2014 5058 2570
rect 800 2008 5058 2014
rect 5122 2008 16189 2576
rect 800 1992 16189 2008
<< via1 >>
rect 222 40051 578 40607
rect 17326 40205 17646 40549
rect 22672 40191 22992 40535
rect 822 39002 1178 39559
rect 17326 39061 17646 39405
rect 22672 39046 22992 39390
rect 14000 36764 14052 36816
rect 14000 36166 14052 36218
rect 2047 34987 2535 35093
rect 222 3619 578 4175
rect 5058 3613 5122 4181
rect 4114 2886 4263 2974
rect 5004 2886 5092 2974
rect 2053 2674 2616 2788
rect 3330 2668 3478 2794
rect 5049 2751 5101 2803
rect 8779 2808 8867 2862
rect 8779 2774 8813 2808
rect 8813 2774 8867 2808
rect 20759 2620 20825 2672
rect 822 2014 1178 2570
rect 5058 2008 5122 2576
<< metal2 >>
rect 21036 44325 21092 44335
rect 14946 43925 15046 43947
rect 14946 43869 14968 43925
rect 15024 43869 15046 43925
rect 20763 43925 20819 43935
rect 200 40607 600 40629
rect 200 40051 222 40607
rect 578 40051 600 40607
rect 200 40029 600 40051
rect 800 39559 1200 39581
rect 800 39002 822 39559
rect 1178 39002 1200 39559
rect 800 38980 1200 39002
rect 13984 36822 14068 36832
rect 13984 36758 13994 36822
rect 14058 36758 14068 36822
rect 13984 36748 14068 36758
rect 2031 36576 3072 36592
rect 2031 36408 2047 36576
rect 3056 36408 3072 36576
rect 13532 36524 13596 36534
rect 13532 36450 13596 36460
rect 2031 35109 3072 36408
rect 13984 36223 14068 36233
rect 13984 36159 13994 36223
rect 14058 36159 14068 36223
rect 13984 36149 14068 36159
rect 2031 35093 3073 35109
rect 2031 34987 2047 35093
rect 2535 34987 2568 35093
rect 2632 34987 3073 35093
rect 2031 34971 3073 34987
rect 2031 34823 2638 34971
rect 2031 30363 2512 34823
rect 2568 30363 2638 34823
rect 222 4175 578 4185
rect 200 3849 222 3945
rect 578 3849 600 3945
rect 222 3609 578 3619
rect 2031 2788 2638 30363
rect 8763 4495 8883 4517
rect 8763 4419 8785 4495
rect 8861 4419 8883 4495
rect 5042 4181 5138 4197
rect 5042 3613 5058 4181
rect 5122 3613 5138 4181
rect 5042 3597 5138 3613
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 8763 2862 8883 4419
rect 14946 4495 15046 43869
rect 17708 43525 17804 43545
rect 17708 43469 17728 43525
rect 17784 43469 17804 43525
rect 17708 43449 17804 43469
rect 17326 40549 17646 40559
rect 17326 40195 17646 40205
rect 17326 39405 17646 39415
rect 17326 39051 17646 39061
rect 17726 36832 17786 43449
rect 20761 39826 20821 43869
rect 17714 36822 17798 36832
rect 17714 36758 17724 36822
rect 17788 36758 17798 36822
rect 17714 36748 17798 36758
rect 14946 4419 14966 4495
rect 15026 4419 15046 4495
rect 14946 4397 15046 4419
rect 2031 2674 2053 2788
rect 2616 2674 2638 2788
rect 2031 2652 2638 2674
rect 3314 2794 3494 2810
rect 3314 2668 3330 2794
rect 3478 2668 3494 2794
rect 5047 2805 5103 2815
rect 5047 2739 5103 2749
rect 8763 2774 8779 2862
rect 8867 2774 8883 2862
rect 3314 2652 3494 2668
rect 800 2576 5138 2592
rect 800 2570 5058 2576
rect 800 2014 822 2570
rect 1178 2014 5058 2570
rect 800 2008 5058 2014
rect 5122 2008 5138 2576
rect 800 1992 5138 2008
rect 8763 1411 8883 2774
rect 20759 2672 20825 39826
rect 21034 39730 21094 44269
rect 23984 43525 24040 43535
rect 22672 40535 22992 40545
rect 22672 40181 22992 40191
rect 23982 39730 24042 43469
rect 21968 36230 22034 39485
rect 22672 39390 22992 39400
rect 22672 39036 22992 39046
rect 21959 36225 22043 36230
rect 21959 36157 21969 36225
rect 22033 36157 22043 36225
rect 21959 36147 22043 36157
rect 20759 2614 20825 2620
rect 8763 1275 8785 1411
rect 8861 1275 8883 1411
rect 8763 1253 8883 1275
<< via2 >>
rect 21036 44269 21092 44325
rect 14968 43869 15024 43925
rect 20763 43869 20819 43925
rect 222 40051 578 40607
rect 822 39002 1178 39559
rect 13994 36816 14058 36822
rect 13994 36764 14000 36816
rect 14000 36764 14052 36816
rect 14052 36764 14058 36816
rect 13994 36758 14058 36764
rect 2047 36408 3056 36576
rect 13532 36460 13596 36524
rect 13994 36218 14058 36223
rect 13994 36166 14000 36218
rect 14000 36166 14052 36218
rect 14052 36166 14058 36218
rect 13994 36159 14058 36166
rect 2568 34987 2632 35093
rect 2512 30363 2568 34823
rect 222 3619 578 4175
rect 8785 4419 8861 4495
rect 5058 3613 5122 4181
rect 4114 2886 4263 2974
rect 5004 2886 5092 2974
rect 17728 43469 17784 43525
rect 17326 40205 17646 40549
rect 17326 39061 17646 39405
rect 17724 36758 17788 36822
rect 14966 4419 15026 4495
rect 3330 2668 3478 2794
rect 5047 2803 5103 2805
rect 5047 2751 5049 2803
rect 5049 2751 5101 2803
rect 5101 2751 5103 2803
rect 5047 2749 5103 2751
rect 822 2014 1178 2570
rect 5058 2008 5122 2576
rect 23984 43469 24040 43525
rect 22672 40191 22992 40535
rect 22672 39046 22992 39390
rect 21969 36157 22033 36225
rect 8785 1275 8861 1411
<< metal3 >>
rect 18810 44345 18910 44347
rect 18810 44341 21115 44345
rect 18810 44253 18816 44341
rect 18904 44325 21115 44341
rect 18904 44269 21036 44325
rect 21092 44269 21115 44325
rect 18904 44253 21115 44269
rect 18810 44249 21115 44253
rect 18810 44247 18910 44249
rect 200 43941 10082 43945
rect 14946 43941 15046 43947
rect 18258 43945 18358 43947
rect 18258 43941 20841 43945
rect 200 43929 6120 43941
rect 200 43864 216 43929
rect 584 43864 6120 43929
rect 200 43853 6120 43864
rect 6208 43853 6672 43941
rect 6760 43853 7224 43941
rect 7312 43853 7776 43941
rect 7864 43853 8328 43941
rect 8416 43853 8880 43941
rect 8968 43853 9432 43941
rect 9520 43853 9984 43941
rect 10072 43853 10082 43941
rect 14942 43853 14952 43941
rect 15040 43853 15050 43941
rect 18258 43853 18264 43941
rect 18352 43925 20841 43941
rect 18352 43869 20763 43925
rect 20819 43869 20841 43925
rect 18352 43853 20841 43869
rect 200 43849 10082 43853
rect 14946 43847 15046 43853
rect 18258 43849 20841 43853
rect 18258 43847 18358 43849
rect 17154 43545 17254 43547
rect 800 43541 17254 43545
rect 800 43529 10536 43541
rect 800 43465 816 43529
rect 1184 43465 10536 43529
rect 800 43453 10536 43465
rect 10624 43453 11088 43541
rect 11176 43453 11640 43541
rect 11728 43453 12192 43541
rect 12280 43453 12744 43541
rect 12832 43453 13296 43541
rect 13384 43453 13848 43541
rect 13936 43453 14400 43541
rect 14488 43453 15504 43541
rect 15592 43453 16056 43541
rect 16144 43453 16608 43541
rect 16696 43453 17160 43541
rect 17248 43453 17254 43541
rect 800 43449 17254 43453
rect 17154 43447 17254 43449
rect 17706 43541 17806 43547
rect 17706 43453 17712 43541
rect 17800 43453 17806 43541
rect 17706 43447 17806 43453
rect 23778 43545 23878 43547
rect 23778 43541 24062 43545
rect 23778 43453 23784 43541
rect 23872 43525 24062 43541
rect 23872 43469 23984 43525
rect 24040 43469 24062 43525
rect 23872 43453 24062 43469
rect 23778 43449 24062 43453
rect 23778 43447 23878 43449
rect 200 40607 24146 40629
rect 200 40051 222 40607
rect 578 40549 24146 40607
rect 578 40205 17326 40549
rect 17646 40535 24146 40549
rect 17646 40205 22672 40535
rect 578 40191 22672 40205
rect 22992 40191 24146 40535
rect 578 40051 24146 40191
rect 200 40029 24146 40051
rect 800 39559 24146 39581
rect 800 39002 822 39559
rect 1178 39405 24146 39559
rect 1178 39061 17326 39405
rect 17646 39390 24146 39405
rect 17646 39061 22672 39390
rect 1178 39046 22672 39061
rect 22992 39046 24146 39390
rect 1178 39002 24146 39046
rect 800 38981 24146 39002
rect 800 38980 1200 38981
rect 200 37465 14366 37487
rect 200 37109 222 37465
rect 578 37109 14366 37465
rect 200 37087 14366 37109
rect 13984 36822 14068 36832
rect 13984 36758 13994 36822
rect 14058 36820 14068 36822
rect 17714 36822 17798 36832
rect 17714 36820 17724 36822
rect 14058 36760 17724 36820
rect 14058 36758 14068 36760
rect 13984 36748 14068 36758
rect 17714 36758 17724 36760
rect 17788 36758 17798 36822
rect 17714 36748 17798 36758
rect 2031 36576 13606 36592
rect 2031 36408 2047 36576
rect 3056 36524 13606 36576
rect 3056 36460 13532 36524
rect 13596 36460 13606 36524
rect 3056 36408 13606 36460
rect 2031 36392 13606 36408
rect 13984 36223 14068 36233
rect 13984 36159 13994 36223
rect 14058 36221 14068 36223
rect 21959 36225 22043 36230
rect 21959 36221 21969 36225
rect 14058 36161 21969 36221
rect 14058 36159 14068 36161
rect 13984 36149 14068 36159
rect 21959 36157 21969 36161
rect 22033 36157 22043 36225
rect 21959 36147 22043 36157
rect 800 35865 14366 35887
rect 800 35509 822 35865
rect 1178 35509 14366 35865
rect 800 35487 14366 35509
rect 2502 34823 2578 34828
rect 2502 30363 2512 34823
rect 2568 30363 2578 34823
rect 2502 30334 2578 30363
rect 8763 4495 15046 4517
rect 8763 4419 8785 4495
rect 8861 4419 14966 4495
rect 15026 4419 15046 4495
rect 8763 4397 15046 4419
rect 200 4181 5138 4197
rect 200 4175 5058 4181
rect 200 3619 222 4175
rect 578 3619 5058 4175
rect 200 3613 5058 3619
rect 5122 3613 5138 4181
rect 200 3597 5138 3613
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 3314 2805 5113 2810
rect 3314 2794 5047 2805
rect 3314 2668 3330 2794
rect 3478 2749 5047 2794
rect 5103 2749 5113 2805
rect 3478 2744 5113 2749
rect 3478 2668 5110 2744
rect 3314 2663 5110 2668
rect 3314 2652 5108 2663
rect 800 2576 5138 2592
rect 800 2570 5058 2576
rect 800 2014 822 2570
rect 1178 2014 5058 2570
rect 800 2008 5058 2014
rect 5122 2008 5138 2576
rect 800 1992 5138 2008
rect 8763 1411 8883 1433
rect 8763 1275 8785 1411
rect 8861 1275 8883 1411
rect 8763 1253 8883 1275
<< via3 >>
rect 18816 44253 18904 44341
rect 216 43864 584 43929
rect 6120 43853 6208 43941
rect 6672 43853 6760 43941
rect 7224 43853 7312 43941
rect 7776 43853 7864 43941
rect 8328 43853 8416 43941
rect 8880 43853 8968 43941
rect 9432 43853 9520 43941
rect 9984 43853 10072 43941
rect 14952 43925 15040 43941
rect 14952 43869 14968 43925
rect 14968 43869 15024 43925
rect 15024 43869 15040 43925
rect 14952 43853 15040 43869
rect 18264 43853 18352 43941
rect 816 43465 1184 43529
rect 10536 43453 10624 43541
rect 11088 43453 11176 43541
rect 11640 43453 11728 43541
rect 12192 43453 12280 43541
rect 12744 43453 12832 43541
rect 13296 43453 13384 43541
rect 13848 43453 13936 43541
rect 14400 43453 14488 43541
rect 15504 43453 15592 43541
rect 16056 43453 16144 43541
rect 16608 43453 16696 43541
rect 17160 43453 17248 43541
rect 17712 43525 17800 43541
rect 17712 43469 17728 43525
rect 17728 43469 17784 43525
rect 17784 43469 17800 43525
rect 17712 43453 17800 43469
rect 23784 43453 23872 43541
rect 222 40051 578 40607
rect 822 39002 1178 39559
rect 222 37109 578 37465
rect 822 35509 1178 35865
rect 222 3619 578 4175
rect 4114 2886 4263 2974
rect 3330 2668 3478 2794
rect 822 2014 1178 2570
rect 8785 1275 8861 1411
<< metal4 >>
rect 200 43929 600 44152
rect 200 43864 216 43929
rect 584 43864 600 43929
rect 200 40607 600 43864
rect 200 40051 222 40607
rect 578 40051 600 40607
rect 200 37465 600 40051
rect 200 37109 222 37465
rect 578 37109 600 37465
rect 200 4175 600 37109
rect 200 3619 222 4175
rect 578 3619 600 4175
rect 200 1000 600 3619
rect 800 43529 1200 44152
rect 6134 43945 6194 45152
rect 6686 43945 6746 45152
rect 7238 43945 7298 45152
rect 7790 43945 7850 45152
rect 8342 43945 8402 45152
rect 8894 43945 8954 45152
rect 9446 43945 9506 45152
rect 9998 43945 10058 45152
rect 6116 43941 6212 43945
rect 6116 43853 6120 43941
rect 6208 43853 6212 43941
rect 6116 43849 6212 43853
rect 6668 43941 6764 43945
rect 6668 43853 6672 43941
rect 6760 43853 6764 43941
rect 6668 43849 6764 43853
rect 7220 43941 7316 43945
rect 7220 43853 7224 43941
rect 7312 43853 7316 43941
rect 7220 43849 7316 43853
rect 7772 43941 7868 43945
rect 7772 43853 7776 43941
rect 7864 43853 7868 43941
rect 7772 43849 7868 43853
rect 8324 43941 8420 43945
rect 8324 43853 8328 43941
rect 8416 43853 8420 43941
rect 8324 43849 8420 43853
rect 8876 43941 8972 43945
rect 8876 43853 8880 43941
rect 8968 43853 8972 43941
rect 8876 43849 8972 43853
rect 9428 43941 9524 43945
rect 9428 43853 9432 43941
rect 9520 43853 9524 43941
rect 9428 43849 9524 43853
rect 9980 43941 10076 43945
rect 9980 43853 9984 43941
rect 10072 43853 10076 43941
rect 9980 43849 10076 43853
rect 10550 43545 10610 45152
rect 11102 43545 11162 45152
rect 11654 43545 11714 45152
rect 12206 43545 12266 45152
rect 12758 43545 12818 45152
rect 13310 43545 13370 45152
rect 13862 43545 13922 45152
rect 14414 43545 14474 45152
rect 14966 43947 15026 45152
rect 14946 43941 15046 43947
rect 14946 43853 14952 43941
rect 15040 43853 15046 43941
rect 14946 43847 15046 43853
rect 15518 43545 15578 45152
rect 16070 43545 16130 45152
rect 16622 43545 16682 45152
rect 17174 43545 17234 45152
rect 17726 43545 17786 45152
rect 18278 43945 18338 45152
rect 18830 44345 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 18812 44341 18908 44345
rect 18812 44253 18816 44341
rect 18904 44253 18908 44341
rect 18812 44249 18908 44253
rect 18260 43941 18356 43945
rect 18260 43853 18264 43941
rect 18352 43853 18356 43941
rect 18260 43849 18356 43853
rect 23798 43545 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 800 43465 816 43529
rect 1184 43465 1200 43529
rect 800 39559 1200 43465
rect 10532 43541 10628 43545
rect 10532 43453 10536 43541
rect 10624 43453 10628 43541
rect 10532 43449 10628 43453
rect 11084 43541 11180 43545
rect 11084 43453 11088 43541
rect 11176 43453 11180 43541
rect 11084 43449 11180 43453
rect 11636 43541 11732 43545
rect 11636 43453 11640 43541
rect 11728 43453 11732 43541
rect 11636 43449 11732 43453
rect 12188 43541 12284 43545
rect 12188 43453 12192 43541
rect 12280 43453 12284 43541
rect 12188 43449 12284 43453
rect 12740 43541 12836 43545
rect 12740 43453 12744 43541
rect 12832 43453 12836 43541
rect 12740 43449 12836 43453
rect 13292 43541 13388 43545
rect 13292 43453 13296 43541
rect 13384 43453 13388 43541
rect 13292 43449 13388 43453
rect 13844 43541 13940 43545
rect 13844 43453 13848 43541
rect 13936 43453 13940 43541
rect 13844 43449 13940 43453
rect 14396 43541 14492 43545
rect 14396 43453 14400 43541
rect 14488 43453 14492 43541
rect 14396 43449 14492 43453
rect 15500 43541 15596 43545
rect 15500 43453 15504 43541
rect 15592 43453 15596 43541
rect 15500 43449 15596 43453
rect 16052 43541 16148 43545
rect 16052 43453 16056 43541
rect 16144 43453 16148 43541
rect 16052 43449 16148 43453
rect 16604 43541 16700 43545
rect 16604 43453 16608 43541
rect 16696 43453 16700 43541
rect 16604 43449 16700 43453
rect 17156 43541 17252 43545
rect 17156 43453 17160 43541
rect 17248 43453 17252 43541
rect 17156 43449 17252 43453
rect 17708 43541 17804 43545
rect 17708 43453 17712 43541
rect 17800 43453 17804 43541
rect 17708 43449 17804 43453
rect 23780 43541 23876 43545
rect 23780 43453 23784 43541
rect 23872 43453 23876 43541
rect 23780 43449 23876 43453
rect 800 39002 822 39559
rect 1178 39002 1200 39559
rect 800 35865 1200 39002
rect 800 35509 822 35865
rect 1178 35509 1200 35865
rect 800 20479 1200 35509
rect 5098 20479 5202 20583
rect 800 19479 10198 20479
rect 800 2570 1200 19479
rect 4099 2974 4279 2990
rect 4099 2886 4114 2974
rect 4263 2886 4279 2974
rect 800 2014 822 2570
rect 1178 2014 1200 2570
rect 800 1000 1200 2014
rect 3314 2794 3494 2810
rect 3314 2668 3330 2794
rect 3478 2668 3494 2794
rect 3314 713 3494 2668
rect 4099 1073 4279 2886
rect 8699 1411 30542 1433
rect 8699 1275 8785 1411
rect 8861 1275 30542 1411
rect 8699 1253 30542 1275
rect 4099 893 26678 1073
rect 3314 533 22814 713
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 533
rect 26498 0 26678 893
rect 30362 0 30542 1253
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 8829 0 1 2544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1715908107
transform 1 0 12693 0 1 2544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1715908107
transform 1 0 16281 0 1 2544
box -38 -48 130 592
use cp7  x1
timestamp 1731242581
transform -1 0 13366 0 1 35787
box -1000 -812 2140 2603
use pfd  x2
timestamp 1731242581
transform -1 0 24092 0 1 39485
box -92 0 6884 640
use vcoB  x3
timestamp 1731242581
transform 1 0 5200 0 1 2294
box -170 55 3759 1652
use sky130_fd_sc_hd__clkinv_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 8921 0 1 2544
box -38 -48 314 592
use lpf  x5
timestamp 1731242581
transform 1 0 2788 0 1 30335
box -240 -9856 9616 5080
use sky130_fd_sc_hd__dfxbp_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 9197 0 1 2544
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  x9
timestamp 1715908107
transform 1 0 10945 0 1 2544
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  x10
timestamp 1715908107
transform 1 0 12785 0 1 2544
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  x11
timestamp 1715908107
transform 1 0 14533 0 1 2544
box -38 -48 1786 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
