magic
tech sky130A
magscale 1 2
timestamp 1731242581
<< error_p >>
rect -367 -856 367 856
<< nwell >>
rect -367 -856 367 856
<< xpolycontact >>
rect 297 424 367 856
rect -367 -856 -297 -424
<< xpolyres >>
rect -367 250 -131 320
rect -367 -424 -297 250
rect -201 -250 -131 250
rect -35 250 201 320
rect -35 -250 35 250
rect -201 -320 35 -250
rect 131 -250 201 250
rect 297 -250 367 424
rect 131 -320 367 -250
<< labels >>
flabel xpolycontact -332 -821 -332 -821 0 FreeSans 80 0 0 0 r0
flabel xpolycontact 332 821 332 821 0 FreeSans 80 0 0 0 r1
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 3.2 m 1 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 100.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
