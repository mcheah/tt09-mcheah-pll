magic
tech sky130A
timestamp 1726261667
<< error_p >>
rect -77 -68 77 68
<< nwell >>
rect -77 -68 77 68
<< scpmoshvt >>
rect -30 -50 30 50
<< pdiff >>
rect -59 -50 -30 50
rect 30 -50 59 50
<< poly >>
rect -30 50 30 63
rect -30 -63 30 -50
<< properties >>
string FIXED_BBOX -101 -133 101 133
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 1.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
