magic
tech sky130A
magscale 1 2
timestamp 1730846090
<< nwell >>
rect -87 -668 87 668
<< xpolycontact >>
rect -35 184 35 616
rect -35 -616 35 -184
<< xpolyres >>
rect -35 -184 35 184
<< viali >>
rect -19 201 19 598
rect -19 -598 19 -201
<< metal1 >>
rect -25 598 25 610
rect -25 201 -19 598
rect 19 201 25 598
rect -25 189 25 201
rect -25 -201 25 -189
rect -25 -598 -19 -201
rect 19 -598 25 -201
rect -25 -610 25 -598
<< labels >>
flabel viali 0 581 0 581 0 FreeSans 80 0 0 0 r0
flabel viali 0 -581 0 -581 0 FreeSans 80 0 0 0 r1
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 12.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
