magic
tech sky130A
magscale 1 2
timestamp 1731242581
<< nwell >>
rect -92 309 6792 630
<< pwell >>
rect -51 69 6753 251
<< locali >>
rect 309 538 374 575
rect 3529 538 3594 575
rect 342 336 374 538
rect 2083 442 2125 458
rect 2108 408 2125 442
rect 2083 269 2125 408
rect 3563 337 3594 538
rect 5303 269 5345 458
rect 6324 303 6656 311
rect 6358 269 6656 303
rect 6324 259 6656 269
<< viali >>
rect 343 575 377 609
rect 3563 575 3597 609
rect 2074 408 2108 442
rect 63 291 97 325
rect 1789 266 1824 301
rect 2188 266 2223 301
rect 2261 266 2296 301
rect 2334 266 2369 301
rect 3012 289 3046 323
rect 3283 291 3317 325
rect 5009 266 5043 300
rect 5502 266 5536 300
rect 5574 266 5608 300
rect 5646 266 5680 300
rect 6324 269 6358 303
rect 6782 263 6816 297
rect 3012 217 3046 251
rect 6706 133 6740 167
<< metal1 >>
rect 38 609 6754 640
rect 38 575 343 609
rect 377 575 3563 609
rect 3597 575 6754 609
rect 38 544 6754 575
rect 2996 482 6825 516
rect 2058 451 2124 458
rect 2058 399 2065 451
rect 2117 399 2124 451
rect 2058 392 2124 399
rect 47 334 113 341
rect 47 282 54 334
rect 106 282 113 334
rect 2996 323 3062 482
rect 5278 451 5344 454
rect 5278 399 5285 451
rect 5337 399 5344 451
rect 5278 392 5344 399
rect 47 275 113 282
rect 1773 301 2385 317
rect 2996 312 3012 323
rect 3046 312 3062 323
rect 3267 334 3333 341
rect 1773 266 1789 301
rect 1824 266 2188 301
rect 2223 266 2261 301
rect 2296 266 2334 301
rect 2369 266 2385 301
rect 1773 250 2385 266
rect 2992 260 3002 312
rect 3056 260 3066 312
rect 3267 282 3274 334
rect 3326 282 3333 334
rect 3267 275 3333 282
rect 4993 300 5696 316
rect 4993 266 5009 300
rect 5043 266 5502 300
rect 5536 266 5574 300
rect 5608 266 5646 300
rect 5680 266 5696 300
rect 2996 251 3062 260
rect 2996 217 3012 251
rect 3046 217 3062 251
rect 4993 250 5696 266
rect 6300 259 6310 311
rect 6362 259 6372 311
rect 6766 297 6825 482
rect 6766 263 6782 297
rect 6816 263 6825 297
rect 6766 251 6825 263
rect 2996 201 3062 217
rect 787 167 917 195
rect 1507 167 1565 195
rect 4007 167 4137 195
rect 4739 167 4785 195
rect 6689 167 6752 183
rect 787 133 6706 167
rect 6740 133 6752 167
rect 787 124 6752 133
rect 38 0 6754 96
<< via1 >>
rect 2065 442 2117 451
rect 2065 408 2074 442
rect 2074 408 2108 442
rect 2108 408 2117 442
rect 2065 399 2117 408
rect 54 325 106 334
rect 54 291 63 325
rect 63 291 97 325
rect 97 291 106 325
rect 54 282 106 291
rect 5285 399 5337 451
rect 3002 289 3012 312
rect 3012 289 3046 312
rect 3046 289 3056 312
rect 3002 260 3056 289
rect 3274 325 3326 334
rect 3274 291 3283 325
rect 3283 291 3317 325
rect 3317 291 3326 325
rect 3274 282 3326 291
rect 6310 303 6362 311
rect 6310 269 6324 303
rect 6324 269 6358 303
rect 6358 269 6362 303
rect 6310 259 6362 269
<< metal2 >>
rect 47 334 113 640
rect 47 282 54 334
rect 106 282 113 334
rect 47 275 113 282
rect 2058 451 2124 458
rect 2058 399 2065 451
rect 2117 399 2124 451
rect 2058 0 2124 399
rect 3002 322 3054 640
rect 5278 451 5344 454
rect 5278 399 5285 451
rect 5337 399 5344 451
rect 3267 334 3333 341
rect 3002 312 3056 322
rect 3002 250 3056 260
rect 3267 282 3274 334
rect 3326 282 3333 334
rect 3267 0 3333 282
rect 5278 0 5344 399
rect 6310 311 6362 640
rect 6310 249 6362 259
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 5374 0 1 48
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1715908107
transform 1 0 -54 0 1 48
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 38 0 1 48
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x2
timestamp 1715908107
transform 1 0 3258 0 1 48
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_8  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 2154 0 1 48
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x4
timestamp 1715908107
transform 1 0 5466 0 1 48
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 6570 0 1 48
box -38 -48 314 592
<< labels >>
flabel metal2 47 574 113 640 0 FreeSans 640 0 0 0 vref
port 0 nsew
flabel metal2 2058 0 2124 66 0 FreeSans 640 0 0 0 upb
flabel metal2 5278 0 5344 66 0 FreeSans 640 0 0 0 downb
port 4 nsew
flabel metal2 6310 588 6362 640 0 FreeSans 320 0 0 0 down
port 5 nsew
flabel metal2 3002 588 3054 640 0 FreeSans 320 0 0 0 up
port 6 nsew
flabel metal2 3267 0 3333 66 0 FreeSans 640 0 0 0 vin
port 2 nsew
flabel metal1 6750 544 6754 640 0 FreeSans 320 0 0 0 vdd
port 7 nsew
flabel metal1 6750 0 6754 96 0 FreeSans 320 0 0 0 vss
port 8 nsew
<< end >>
