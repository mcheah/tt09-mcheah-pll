magic
tech sky130A
magscale 1 2
timestamp 1729864714
<< nwell >>
rect -154 -242 154 242
<< pmos >>
rect -60 -180 60 180
<< pdiff >>
rect -118 168 -60 180
rect -118 -168 -106 168
rect -72 -168 -60 168
rect -118 -180 -60 -168
rect 60 168 118 180
rect 60 -168 72 168
rect 106 -168 118 168
rect 60 -180 118 -168
<< pdiffc >>
rect -106 -168 -72 168
rect 72 -168 106 168
<< poly >>
rect -60 180 60 206
rect -60 -206 60 -180
<< locali >>
rect -106 168 -72 184
rect -106 -184 -72 -168
rect 72 168 106 184
rect 72 -184 106 -168
<< labels >>
flabel pdiffc -89 0 -89 0 0 FreeSans 80 0 0 0 d
flabel pdiffc 89 0 89 0 0 FreeSans 80 0 0 0 s
flabel pmos -60 -180 60 180 0 FreeSans 80 0 0 0 g
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.8 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
