magic
tech sky130A
magscale 1 2
timestamp 1729864714
<< nwell >>
rect -109 -122 109 122
<< pmos >>
rect -15 -60 15 60
<< pdiff >>
rect -73 48 -15 60
rect -73 -48 -61 48
rect -27 -48 -15 48
rect -73 -60 -15 -48
rect 15 48 73 60
rect 15 -48 27 48
rect 61 -48 73 48
rect 15 -60 73 -48
<< pdiffc >>
rect -61 -48 -27 48
rect 27 -48 61 48
<< poly >>
rect -15 60 15 86
rect -15 -86 15 -60
<< locali >>
rect -61 48 -27 64
rect -61 -64 -27 -48
rect 27 48 61 64
rect 27 -64 61 -48
<< labels >>
flabel pdiffc -44 0 -44 0 0 FreeSans 80 0 0 0 d
flabel pdiffc 44 0 44 0 0 FreeSans 80 0 0 0 s
flabel pmos -15 -60 15 60 0 FreeSans 80 0 0 0 g
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.6 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
