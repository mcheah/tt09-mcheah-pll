magic
tech sky130A
magscale 1 2
timestamp 1726197802
<< xpolycontact >>
rect 297 454 367 886
rect -367 -886 -297 -454
<< xpolyres >>
rect -367 280 -131 350
rect -367 -454 -297 280
rect -201 -280 -131 280
rect -35 280 201 350
rect -35 -280 35 280
rect -201 -350 35 -280
rect 131 -280 201 280
rect 297 -280 367 454
rect 131 -350 367 -280
<< labels >>
flabel locali 297 454 367 886 0 FreeSans 160 0 0 0 r0
flabel locali -367 -886 -297 -454 0 FreeSans 160 0 0 0 r1
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 3.5 m 1 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 109.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
