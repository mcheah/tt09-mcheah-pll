magic
tech sky130A
magscale 1 2
timestamp 1726197802
<< nmos >>
rect -60 -50 60 50
<< ndiff >>
rect -118 38 -60 50
rect -118 -38 -106 38
rect -72 -38 -60 38
rect -118 -50 -60 -38
rect 60 38 118 50
rect 60 -38 72 38
rect 106 -38 118 38
rect 60 -50 118 -38
<< ndiffc >>
rect -106 -38 -72 38
rect 72 -38 106 38
<< poly >>
rect -60 50 60 76
rect -60 -76 60 -50
<< locali >>
rect -106 38 -72 54
rect -106 -54 -72 -38
rect 72 38 106 54
rect 72 -54 106 -38
<< labels >>
flabel locali -89 0 -89 0 0 FreeSans 80 0 0 0 d
port 0 nsew
flabel locali 89 0 89 0 0 FreeSans 80 0 0 0 s
port 1 nsew
flabel poly -60 -50 60 50 0 FreeSans 80 0 0 0 g
port 2 nsew
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w .5 l .6 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
