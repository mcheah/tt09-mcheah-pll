magic
tech sky130A
magscale 1 2
timestamp 1726261667
<< error_s >>
rect -218 -415 -160 -285
rect -40 -415 18 -285
rect -313 -837 110 -499
<< nwell >>
rect -313 -837 110 -499
<< pwell >>
rect 10 -259 44 -221
rect -244 -441 44 -259
<< ndiffc >>
rect -210 -333 -176 -299
rect -24 -333 10 -299
rect -210 -401 -176 -367
rect -24 -401 10 -367
<< pdiffc >>
rect -210 -584 -176 -550
rect -24 -584 10 -550
rect -210 -652 -176 -618
rect -24 -652 10 -618
rect -210 -720 -176 -686
rect -24 -720 10 -686
<< poly >>
rect -160 -454 -40 -441
rect -160 -488 -110 -454
rect -76 -488 -40 -454
rect -160 -509 -40 -488
<< polycont >>
rect -110 -488 -76 -454
<< locali >>
rect -292 -255 -209 -221
rect -175 -255 -117 -221
rect -83 -255 -25 -221
rect 9 -255 89 -221
rect -226 -299 -160 -289
rect -226 -333 -210 -299
rect -176 -333 -160 -299
rect -226 -367 -160 -333
rect -226 -401 -210 -367
rect -176 -401 -160 -367
rect -226 -415 -160 -401
rect -24 -299 22 -255
rect 10 -333 22 -299
rect -24 -367 22 -333
rect 10 -401 22 -367
rect -226 -535 -180 -415
rect -24 -417 22 -401
rect -126 -452 -60 -441
rect -126 -454 22 -452
rect -126 -488 -110 -454
rect -76 -488 22 -454
rect -126 -499 22 -488
rect -126 -509 -60 -499
rect -226 -550 -160 -535
rect -226 -584 -210 -550
rect -176 -584 -160 -550
rect -226 -618 -160 -584
rect -226 -652 -210 -618
rect -176 -652 -160 -618
rect -226 -686 -160 -652
rect -226 -720 -210 -686
rect -176 -720 -160 -686
rect -226 -729 -160 -720
rect -24 -550 23 -534
rect 10 -584 23 -550
rect -24 -618 23 -584
rect 10 -652 23 -618
rect -24 -686 23 -652
rect 10 -720 23 -686
rect -24 -765 23 -720
rect -292 -799 -209 -765
rect -175 -799 -117 -765
rect -83 -799 -25 -765
rect 9 -799 89 -765
<< viali >>
rect -209 -255 -175 -221
rect -117 -255 -83 -221
rect -25 -255 9 -221
rect -209 -799 -175 -765
rect -117 -799 -83 -765
rect -25 -799 9 -765
<< metal1 >>
rect -292 -221 89 -190
rect -292 -255 -209 -221
rect -175 -255 -117 -221
rect -83 -255 -25 -221
rect 9 -255 89 -221
rect -292 -286 89 -255
rect -292 -765 89 -734
rect -292 -799 -209 -765
rect -175 -799 -117 -765
rect -83 -799 -25 -765
rect 9 -799 89 -765
rect -292 -830 89 -799
use sky130_fd_pr__nfet_01v8_RFBLNB  XM1
timestamp 1725317697
transform 1 0 -100 0 1 -350
box -118 -91 118 91
use sky130_fd_pr__pfet_01v8_hvt_XPYSBA  XM2
timestamp 1726261667
transform 1 0 -100 0 1 -635
box -154 -136 154 136
<< labels >>
flabel metal1 -292 -286 89 -190 7 FreeSans 360 0 0 0 VSS
port 0 w
flabel metal1 -292 -830 89 -734 7 FreeSans 360 0 0 0 VDD
port 1 w
flabel locali -25 -499 22 -452 3 FreeSans 360 0 0 0 A
port 2 e
flabel locali -226 -499 -180 -452 7 FreeSans 360 0 0 0 Y
port 3 w
flabel pwell 10 -255 44 -221 0 FreeSans 160 0 0 0 VNB
port 4 nsew
flabel nwell 10 -799 44 -765 0 FreeSans 160 0 0 0 VPB
port 5 nsew
<< end >>
