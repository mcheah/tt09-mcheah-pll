magic
tech sky130A
magscale 1 2
timestamp 1729864714
<< nwell >>
rect -154 -152 154 152
<< pmos >>
rect -60 -90 60 90
<< pdiff >>
rect -118 78 -60 90
rect -118 -78 -106 78
rect -72 -78 -60 78
rect -118 -90 -60 -78
rect 60 78 118 90
rect 60 -78 72 78
rect 106 -78 118 78
rect 60 -90 118 -78
<< pdiffc >>
rect -106 -78 -72 78
rect 72 -78 106 78
<< poly >>
rect -60 90 60 116
rect -60 -116 60 -90
<< locali >>
rect -106 78 -72 94
rect -106 -94 -72 -78
rect 72 78 106 94
rect 72 -94 106 -78
<< labels >>
flabel pdiffc -89 0 -89 0 0 FreeSans 80 0 0 0 d
flabel pdiffc 89 0 89 0 0 FreeSans 80 0 0 0 s
flabel pmos -60 -90 60 90 0 FreeSans 80 0 0 0 g
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.9 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
