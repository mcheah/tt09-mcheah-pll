magic
tech sky130A
magscale 1 2
timestamp 1730848472
<< pwell >>
rect -121 -2503 121 2503
<< xpolycontact >>
rect -69 2019 69 2451
rect -69 -2451 69 -2019
<< ppolyres >>
rect -69 -2019 69 2019
<< viali >>
rect -53 2036 53 2433
rect -53 -2433 53 -2036
<< metal1 >>
rect -59 2433 59 2445
rect -59 2036 -53 2433
rect 53 2036 59 2433
rect -59 2024 59 2036
rect -59 -2036 59 -2024
rect -59 -2433 -53 -2036
rect 53 -2433 59 -2036
rect -59 -2445 59 -2433
<< labels >>
flabel viali 0 2416 0 2416 0 FreeSans 80 0 0 0 r0
flabel viali 0 -2416 0 -2416 0 FreeSans 80 0 0 0 r1
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 20.35 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 9.996k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
