magic
tech sky130A
magscale 1 2
timestamp 1726339549
<< metal1 >>
rect 200 3929 5138 3945
rect 200 3865 216 3929
rect 584 3865 5058 3929
rect 5122 3865 5138 3929
rect 200 3849 5138 3865
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 8763 2862 18950 2878
rect 3314 2794 5108 2810
rect 3314 2668 3330 2794
rect 3478 2668 4966 2794
rect 5092 2668 5108 2794
rect 8763 2774 8779 2862
rect 8867 2774 14862 2862
rect 15010 2774 18786 2862
rect 18934 2774 18950 2862
rect 8763 2758 18950 2774
rect 3314 2652 5108 2668
rect 800 2576 5138 2592
rect 800 2512 816 2576
rect 1184 2512 5058 2576
rect 5122 2512 5138 2576
rect 800 2496 5138 2512
<< via1 >>
rect 216 3865 584 3929
rect 5058 3865 5122 3929
rect 4114 2886 4263 2974
rect 5004 2886 5092 2974
rect 3330 2668 3478 2794
rect 4966 2668 5092 2794
rect 8779 2774 8867 2862
rect 14862 2774 15010 2862
rect 18786 2774 18934 2862
rect 816 2512 1184 2576
rect 5058 2512 5122 2576
<< metal2 >>
rect 200 3929 5138 3945
rect 200 3865 216 3929
rect 584 3865 5058 3929
rect 5122 3865 5138 3929
rect 200 3849 5138 3865
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 8763 2862 18950 2878
rect 3314 2794 5108 2810
rect 3314 2668 3330 2794
rect 3478 2668 4966 2794
rect 5092 2668 5108 2794
rect 8763 2774 8779 2862
rect 8867 2774 14862 2862
rect 15010 2774 18786 2862
rect 18934 2774 18950 2862
rect 8763 2758 18950 2774
rect 3314 2652 5108 2668
rect 800 2576 5138 2592
rect 800 2512 816 2576
rect 1184 2512 5058 2576
rect 5122 2512 5138 2576
rect 800 2496 5138 2512
<< via2 >>
rect 216 3865 584 3929
rect 5058 3865 5122 3929
rect 4114 2886 4263 2974
rect 5004 2886 5092 2974
rect 3330 2668 3478 2794
rect 4966 2668 5092 2794
rect 8779 2774 8867 2862
rect 14862 2774 15010 2862
rect 18786 2774 18934 2862
rect 816 2512 1184 2576
rect 5058 2512 5122 2576
<< metal3 >>
rect 200 43941 10082 43945
rect 200 43929 6120 43941
rect 200 43864 216 43929
rect 584 43864 6120 43929
rect 200 43853 6120 43864
rect 6208 43853 6672 43941
rect 6760 43853 7224 43941
rect 7312 43853 7776 43941
rect 7864 43853 8328 43941
rect 8416 43853 8880 43941
rect 8968 43853 9432 43941
rect 9520 43853 9984 43941
rect 10072 43853 10082 43941
rect 200 43849 10082 43853
rect 800 43541 18925 43545
rect 800 43529 10536 43541
rect 800 43465 816 43529
rect 1184 43465 10536 43529
rect 800 43453 10536 43465
rect 10624 43453 11088 43541
rect 11176 43453 11640 43541
rect 11728 43453 12192 43541
rect 12280 43453 12744 43541
rect 12832 43453 13296 43541
rect 13384 43453 13848 43541
rect 13936 43453 14400 43541
rect 14488 43453 15504 43541
rect 15592 43453 16056 43541
rect 16144 43453 16608 43541
rect 16696 43453 17160 43541
rect 17248 43453 17712 43541
rect 17800 43453 18264 43541
rect 18352 43453 18816 43541
rect 18904 43453 18925 43541
rect 800 43449 18925 43453
rect 200 3929 5138 3945
rect 200 3865 216 3929
rect 584 3865 5058 3929
rect 5122 3865 5138 3929
rect 200 3849 5138 3865
rect 4099 2974 5108 2990
rect 4099 2886 4114 2974
rect 4263 2886 5004 2974
rect 5092 2886 5108 2974
rect 4099 2870 5108 2886
rect 8763 2862 18950 2878
rect 3314 2794 5108 2810
rect 3314 2668 3330 2794
rect 3478 2668 4966 2794
rect 5092 2668 5108 2794
rect 8763 2774 8779 2862
rect 8867 2774 14862 2862
rect 15010 2774 18786 2862
rect 18934 2774 18950 2862
rect 8763 2758 18950 2774
rect 3314 2652 5108 2668
rect 800 2576 5138 2592
rect 800 2512 816 2576
rect 1184 2512 5058 2576
rect 5122 2512 5138 2576
rect 800 2496 5138 2512
<< via3 >>
rect 216 43864 584 43929
rect 6120 43853 6208 43941
rect 6672 43853 6760 43941
rect 7224 43853 7312 43941
rect 7776 43853 7864 43941
rect 8328 43853 8416 43941
rect 8880 43853 8968 43941
rect 9432 43853 9520 43941
rect 9984 43853 10072 43941
rect 816 43465 1184 43529
rect 10536 43453 10624 43541
rect 11088 43453 11176 43541
rect 11640 43453 11728 43541
rect 12192 43453 12280 43541
rect 12744 43453 12832 43541
rect 13296 43453 13384 43541
rect 13848 43453 13936 43541
rect 14400 43453 14488 43541
rect 15504 43453 15592 43541
rect 16056 43453 16144 43541
rect 16608 43453 16696 43541
rect 17160 43453 17248 43541
rect 17712 43453 17800 43541
rect 18264 43453 18352 43541
rect 18816 43453 18904 43541
rect 216 3865 584 3929
rect 4114 2886 4263 2974
rect 3330 2668 3478 2794
rect 14862 2774 15010 2862
rect 18786 2774 18934 2862
rect 816 2512 1184 2576
<< metal4 >>
rect 200 43929 600 44152
rect 200 43864 216 43929
rect 584 43864 600 43929
rect 200 3929 600 43864
rect 200 3865 216 3929
rect 584 3865 600 3929
rect 200 1000 600 3865
rect 800 43529 1200 44152
rect 6134 43945 6194 45152
rect 6686 43945 6746 45152
rect 7238 43945 7298 45152
rect 7790 43945 7850 45152
rect 8342 43945 8402 45152
rect 8894 43945 8954 45152
rect 9446 43945 9506 45152
rect 9998 43945 10058 45152
rect 6116 43941 6212 43945
rect 6116 43853 6120 43941
rect 6208 43853 6212 43941
rect 6116 43849 6212 43853
rect 6668 43941 6764 43945
rect 6668 43853 6672 43941
rect 6760 43853 6764 43941
rect 6668 43849 6764 43853
rect 7220 43941 7316 43945
rect 7220 43853 7224 43941
rect 7312 43853 7316 43941
rect 7220 43849 7316 43853
rect 7772 43941 7868 43945
rect 7772 43853 7776 43941
rect 7864 43853 7868 43941
rect 7772 43849 7868 43853
rect 8324 43941 8420 43945
rect 8324 43853 8328 43941
rect 8416 43853 8420 43941
rect 8324 43849 8420 43853
rect 8876 43941 8972 43945
rect 8876 43853 8880 43941
rect 8968 43853 8972 43941
rect 8876 43849 8972 43853
rect 9428 43941 9524 43945
rect 9428 43853 9432 43941
rect 9520 43853 9524 43941
rect 9428 43849 9524 43853
rect 9980 43941 10076 43945
rect 9980 43853 9984 43941
rect 10072 43853 10076 43941
rect 9980 43849 10076 43853
rect 10550 43545 10610 45152
rect 11102 43545 11162 45152
rect 11654 43545 11714 45152
rect 12206 43545 12266 45152
rect 12758 43545 12818 45152
rect 13310 43545 13370 45152
rect 13862 43545 13922 45152
rect 14414 43545 14474 45152
rect 800 43465 816 43529
rect 1184 43465 1200 43529
rect 800 2576 1200 43465
rect 10532 43541 10628 43545
rect 10532 43453 10536 43541
rect 10624 43453 10628 43541
rect 10532 43449 10628 43453
rect 11084 43541 11180 43545
rect 11084 43453 11088 43541
rect 11176 43453 11180 43541
rect 11084 43449 11180 43453
rect 11636 43541 11732 43545
rect 11636 43453 11640 43541
rect 11728 43453 11732 43541
rect 11636 43449 11732 43453
rect 12188 43541 12284 43545
rect 12188 43453 12192 43541
rect 12280 43453 12284 43541
rect 12188 43449 12284 43453
rect 12740 43541 12836 43545
rect 12740 43453 12744 43541
rect 12832 43453 12836 43541
rect 12740 43449 12836 43453
rect 13292 43541 13388 43545
rect 13292 43453 13296 43541
rect 13384 43453 13388 43541
rect 13292 43449 13388 43453
rect 13844 43541 13940 43545
rect 13844 43453 13848 43541
rect 13936 43453 13940 43541
rect 13844 43449 13940 43453
rect 14396 43541 14492 43545
rect 14396 43453 14400 43541
rect 14488 43453 14492 43541
rect 14396 43449 14492 43453
rect 4099 2974 4279 2990
rect 4099 2886 4114 2974
rect 4263 2886 4279 2974
rect 800 2512 816 2576
rect 1184 2512 1200 2576
rect 800 1000 1200 2512
rect 3314 2794 3494 2810
rect 3314 2668 3330 2794
rect 3478 2668 3494 2794
rect 3314 713 3494 2668
rect 4099 1073 4279 2886
rect 14966 2878 15026 45152
rect 15518 43545 15578 45152
rect 16070 43545 16130 45152
rect 16622 43545 16682 45152
rect 17174 43545 17234 45152
rect 17726 43545 17786 45152
rect 18278 43545 18338 45152
rect 18830 43545 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 15500 43541 15596 43545
rect 15500 43453 15504 43541
rect 15592 43453 15596 43541
rect 15500 43449 15596 43453
rect 16052 43541 16148 43545
rect 16052 43453 16056 43541
rect 16144 43453 16148 43541
rect 16052 43449 16148 43453
rect 16604 43541 16700 43545
rect 16604 43453 16608 43541
rect 16696 43453 16700 43541
rect 16604 43449 16700 43453
rect 17156 43541 17252 43545
rect 17156 43453 17160 43541
rect 17248 43453 17252 43541
rect 17156 43449 17252 43453
rect 17708 43541 17804 43545
rect 17708 43453 17712 43541
rect 17800 43453 17804 43541
rect 17708 43449 17804 43453
rect 18260 43541 18356 43545
rect 18260 43453 18264 43541
rect 18352 43453 18356 43541
rect 18260 43449 18356 43453
rect 18812 43541 18908 43545
rect 18812 43453 18816 43541
rect 18904 43453 18908 43541
rect 18812 43449 18908 43453
rect 14846 2862 15026 2878
rect 14846 2774 14862 2862
rect 15010 2774 15026 2862
rect 14846 2758 15026 2774
rect 18770 2862 18950 2878
rect 18770 2774 18786 2862
rect 18934 2774 18950 2862
rect 4099 893 15086 1073
rect 3314 533 11222 713
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 533
rect 14906 0 15086 893
rect 18770 0 18950 2774
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use vcoB  vcoB_0
timestamp 1726339549
transform 1 0 5200 0 1 2294
box -170 55 3759 1652
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
