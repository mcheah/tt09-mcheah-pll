magic
tech sky130A
magscale 1 2
timestamp 1731242581
<< error_s >>
rect -902 1603 434 1777
rect -234 998 608 1482
rect -168 564 318 744
rect -168 260 608 564
rect -20 -755 38 -665
rect 338 -755 396 -665
rect 507 -836 541 -802
rect -198 -1243 -140 -883
rect -20 -1243 38 -883
rect 158 -1243 216 -883
<< poly >>
rect -140 1040 -20 1446
rect 38 1040 158 1446
rect 216 1040 336 1446
rect 394 1040 514 1446
rect -140 933 514 1040
rect -140 909 -31 933
rect -74 899 -31 909
rect 3 909 147 933
rect 3 899 46 909
rect -74 296 46 899
rect 104 899 147 909
rect 181 909 514 933
rect 181 899 224 909
rect 104 322 224 899
rect 394 248 514 502
rect 394 214 437 248
rect 471 214 514 248
rect 394 198 514 214
rect 38 -583 338 -567
rect 38 -617 171 -583
rect 205 -617 338 -583
rect 38 -781 338 -617
rect -140 -1269 -20 -883
rect 38 -1269 158 -883
rect -140 -1291 158 -1269
rect -140 -1325 -97 -1291
rect -63 -1325 81 -1291
rect 115 -1325 158 -1291
rect -140 -1341 158 -1325
<< polycont >>
rect -31 899 3 933
rect 147 899 181 933
rect 437 214 471 248
rect 171 -617 205 -583
rect -97 -1325 -63 -1291
rect 81 -1325 115 -1291
<< locali >>
rect -50 1655 382 1725
rect -8 1474 382 1655
rect -186 1017 -152 1424
rect -8 1056 26 1474
rect 170 1017 204 1424
rect 348 1056 382 1474
rect 526 1033 560 1424
rect 510 1017 576 1033
rect -186 983 526 1017
rect 560 983 576 1017
rect 510 967 576 983
rect -47 933 19 949
rect 131 933 197 949
rect -188 899 -31 933
rect 3 899 147 933
rect 181 899 270 933
rect -188 796 -154 899
rect -47 883 19 899
rect 131 883 197 899
rect -204 780 -138 796
rect -204 746 -188 780
rect -154 746 -138 780
rect -204 730 -138 746
rect -120 248 -86 686
rect 58 334 92 670
rect 236 506 270 899
rect 236 318 382 506
rect 526 334 560 967
rect 421 248 487 264
rect -120 214 437 248
rect 471 214 487 248
rect 421 198 487 214
rect -204 -545 -138 -529
rect -204 -579 -188 -545
rect -154 -579 -138 -545
rect -204 -595 -138 -579
rect 155 -583 221 -567
rect -186 -1247 -152 -595
rect 155 -617 171 -583
rect 205 -617 384 -583
rect 155 -633 221 -617
rect -8 -1247 26 -661
rect 350 -759 384 -617
rect -113 -1291 -47 -1275
rect 65 -1291 131 -1275
rect 170 -1291 204 -895
rect -113 -1325 -97 -1291
rect -63 -1325 81 -1291
rect 115 -1325 526 -1291
rect -113 -1341 -47 -1325
rect 65 -1341 131 -1325
<< viali >>
rect 526 983 560 1017
rect -188 746 -154 780
rect 437 214 471 248
rect -188 -579 -154 -545
rect 171 -617 205 -583
rect 526 -1325 560 -1291
<< metal1 >>
rect -850 1671 -816 1705
rect 510 1026 576 1033
rect 507 974 517 1026
rect 569 974 579 1026
rect 510 967 576 974
rect -207 789 -135 796
rect -207 737 -197 789
rect -145 737 -135 789
rect -204 730 -138 737
rect 418 205 428 257
rect 480 205 490 257
rect -204 -536 -138 -529
rect -207 -588 -197 -536
rect -145 -588 -135 -536
rect 155 -574 221 -567
rect -204 -595 -138 -588
rect 152 -626 162 -574
rect 214 -626 224 -574
rect 155 -633 221 -626
rect 507 -836 541 -802
rect 507 -1334 517 -1282
rect 569 -1334 579 -1282
<< via1 >>
rect 517 1017 569 1026
rect 517 983 526 1017
rect 526 983 560 1017
rect 560 983 569 1017
rect 517 974 569 983
rect -197 780 -145 789
rect -197 746 -188 780
rect -188 746 -154 780
rect -154 746 -145 780
rect -197 737 -145 746
rect 428 248 480 257
rect 428 214 437 248
rect 437 214 471 248
rect 471 214 480 248
rect 428 205 480 214
rect -197 -545 -145 -536
rect -197 -579 -188 -545
rect -188 -579 -154 -545
rect -154 -579 -145 -545
rect -197 -588 -145 -579
rect 162 -583 214 -574
rect 162 -617 171 -583
rect 171 -617 205 -583
rect 205 -617 214 -583
rect 162 -626 214 -617
rect 517 -1291 569 -1282
rect 517 -1325 526 -1291
rect 526 -1325 560 -1291
rect 560 -1325 569 -1291
rect 517 -1334 569 -1325
<< metal2 >>
rect 517 1026 569 1036
rect 517 964 569 974
rect -197 789 -145 799
rect -197 727 -145 737
rect -188 -526 -154 727
rect 428 257 480 267
rect 171 214 428 248
rect -197 -536 -145 -526
rect 171 -564 205 214
rect 428 195 480 205
rect -197 -598 -145 -588
rect 162 -574 214 -564
rect 162 -636 214 -626
rect 526 -1272 560 964
rect 517 -1282 569 -1272
rect 517 -1344 569 -1334
use sky130_fd_pr__nfet_01v8_ZJWC73  XM1
timestamp 1729864714
transform 1 0 -80 0 1 -1063
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_ZJWC73  XM2
timestamp 1729864714
transform -1 0 98 0 1 -1063
box -118 -206 118 206
use sky130_fd_pr__pfet_01v8_AH2TBC  XM3
timestamp 1729864714
transform -1 0 164 0 1 502
box -154 -242 154 242
use sky130_fd_pr__pfet_01v8_AH6ZBC  XM4
timestamp 1730210991
transform 1 0 187 0 1 1240
box -421 -242 421 242
use sky130_fd_pr__pfet_01v8_AH2TBC  XM5
timestamp 1729864714
transform 1 0 -14 0 -1 502
box -154 -242 154 242
use sky130_fd_pr__nfet_01v8_HE5L4J  XM6
timestamp 1729864714
transform -1 0 188 0 1 -710
box -208 -71 208 71
use sky130_fd_pr__pfet_01v8_EP2VBC  XM7
timestamp 1729864714
transform -1 0 454 0 1 412
box -154 -152 154 152
use sky130_fd_pr__res_xhigh_po_0p35_QBQWER  XR1 $PDKPATH/libs.tech/magic
timestamp 1730846090
transform 0 1 -234 -1 0 1690
box -87 -668 87 668
<< labels >>
flabel metal1 -850 1671 -816 1705 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 -193 770 -159 771 0 FreeSans 256 0 0 0 vpb
port 2 nsew
flabel locali -8 -710 26 -676 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 507 -836 541 -802 0 FreeSans 240 0 0 0 vnb
port 4 nsew
<< end >>
