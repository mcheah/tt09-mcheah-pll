magic
tech sky130A
magscale 1 2
timestamp 1731242581
<< nwell >>
rect -546 709 1649 2603
<< pwell >>
rect -553 -812 1619 701
<< psubdiff >>
rect -517 631 -421 665
rect 1487 631 1583 665
rect -517 569 -483 631
rect 1549 569 1583 631
rect -517 -742 -483 -680
rect 1549 -742 1583 -680
rect -517 -776 -421 -742
rect 1487 -776 1583 -742
<< nsubdiff >>
rect -510 2533 -414 2567
rect 1517 2533 1613 2567
rect -510 2471 -476 2533
rect 1579 2471 1613 2533
rect -510 779 -476 841
rect 1579 779 1613 841
rect -510 745 -414 779
rect 1517 745 1613 779
<< psubdiffcont >>
rect -421 631 1487 665
rect -517 -680 -483 569
rect 1549 -680 1583 569
rect -421 -776 1487 -742
<< nsubdiffcont >>
rect -414 2533 1517 2567
rect -510 841 -476 2471
rect 1579 841 1613 2471
rect -414 745 1517 779
<< poly >>
rect 59 2145 179 2156
rect 59 2111 102 2145
rect 136 2111 179 2145
rect -119 1615 1 2048
rect -119 1581 -76 1615
rect -42 1581 1 1615
rect -319 1036 -289 1196
rect -337 1020 -271 1036
rect -337 986 -321 1020
rect -287 986 -271 1020
rect -337 970 -271 986
rect -119 930 1 1581
rect 59 1615 179 2111
rect 59 1581 102 1615
rect 136 1581 179 1615
rect 59 1549 179 1581
rect 74 1429 179 1549
rect 59 1397 179 1429
rect 59 1363 102 1397
rect 136 1363 179 1397
rect 59 930 179 1363
rect 237 1615 357 2048
rect 237 1581 280 1615
rect 314 1581 357 1615
rect 237 1397 357 1581
rect 237 1363 280 1397
rect 314 1363 357 1397
rect 237 956 357 1363
rect -119 563 1 579
rect -119 529 -76 563
rect -42 529 1 563
rect -335 421 -269 437
rect -335 387 -319 421
rect -285 387 -269 421
rect -335 371 -269 387
rect -319 243 -289 371
rect -119 -169 1 529
rect 59 49 179 482
rect 59 15 102 49
rect 136 15 179 49
rect 59 -17 179 15
rect 74 -137 179 -17
rect -119 -203 -76 -169
rect -42 -203 1 -169
rect -119 -636 1 -203
rect 59 -169 179 -137
rect 59 -203 102 -169
rect 136 -203 179 -169
rect 59 -657 179 -203
rect 237 49 357 482
rect 237 15 280 49
rect 314 15 357 49
rect 237 -169 357 15
rect 237 -203 280 -169
rect 314 -203 357 -169
rect 237 -610 357 -203
rect 59 -691 102 -657
rect 136 -691 179 -657
rect 59 -731 179 -691
<< polycont >>
rect 102 2111 136 2145
rect -76 1581 -42 1615
rect -321 986 -287 1020
rect 102 1581 136 1615
rect 102 1363 136 1397
rect 280 1581 314 1615
rect 280 1363 314 1397
rect -76 529 -42 563
rect -319 387 -285 421
rect 102 15 136 49
rect -76 -203 -42 -169
rect 102 -203 136 -169
rect 280 15 314 49
rect 280 -203 314 -169
rect 102 -691 136 -657
<< locali >>
rect -510 2533 -414 2567
rect 1517 2533 1613 2567
rect -510 2471 -476 2533
rect 162 2473 178 2533
rect 238 2473 254 2533
rect 162 2457 254 2473
rect 1579 2471 1613 2533
rect 86 2146 152 2161
rect 86 2145 573 2146
rect -165 2111 102 2145
rect 136 2111 573 2145
rect -165 1700 -131 2111
rect 86 2095 152 2111
rect 13 1700 47 2036
rect -92 1615 -26 1631
rect -476 1570 -400 1586
rect -416 1510 -400 1570
rect -476 1494 -400 1510
rect -165 1581 -76 1615
rect -42 1581 -26 1615
rect -165 1456 -131 1581
rect -92 1565 -26 1581
rect 86 1615 152 1631
rect 86 1581 102 1615
rect 136 1581 152 1615
rect 86 1565 152 1581
rect 13 1506 47 1522
rect 191 1521 225 2036
rect 369 1885 403 2036
rect 473 1901 539 1917
rect 473 1885 489 1901
rect 369 1867 489 1885
rect 523 1867 539 1901
rect 369 1851 539 1867
rect 369 1700 403 1851
rect 264 1615 330 1631
rect 264 1581 280 1615
rect 314 1581 330 1615
rect 264 1565 330 1581
rect 405 1615 471 1631
rect 405 1581 421 1615
rect 455 1581 471 1615
rect 405 1565 471 1581
rect 175 1506 241 1521
rect 13 1505 241 1506
rect 13 1472 191 1505
rect 13 1456 47 1472
rect 175 1471 191 1472
rect 225 1471 241 1505
rect 175 1455 241 1471
rect -442 1397 -376 1413
rect 86 1397 152 1413
rect -442 1363 -426 1397
rect -392 1363 47 1397
rect -442 1347 -376 1363
rect -265 1313 -199 1329
rect -365 1281 -299 1297
rect -365 1247 -349 1281
rect -315 1247 -299 1281
rect -365 1231 -299 1247
rect -265 1279 -249 1313
rect -215 1279 -199 1313
rect -265 1263 -199 1279
rect -365 1088 -331 1231
rect -265 1072 -222 1263
rect -337 1020 -271 1036
rect -337 986 -321 1020
rect -287 986 -271 1020
rect -165 1018 -131 1304
rect -337 970 -271 986
rect -231 1002 -131 1018
rect -231 968 -215 1002
rect -181 968 -131 1002
rect 13 968 47 1363
rect 86 1363 102 1397
rect 136 1363 152 1397
rect 86 1347 152 1363
rect 191 968 225 1455
rect 280 1413 314 1565
rect 1547 1560 1579 1576
rect 981 1423 1047 1439
rect 264 1397 330 1413
rect 264 1363 280 1397
rect 314 1363 330 1397
rect 981 1389 997 1423
rect 1031 1389 1047 1423
rect 981 1373 1047 1389
rect 264 1347 330 1363
rect -231 952 -131 968
rect -510 779 -476 841
rect -92 863 -26 879
rect 369 863 403 1320
rect 997 1319 1031 1373
rect 1547 1360 1563 1560
rect 1547 1344 1579 1360
rect -92 829 -76 863
rect -42 829 403 863
rect -92 813 -26 829
rect 1579 779 1613 841
rect -510 745 -414 779
rect 1517 745 1613 779
rect -517 631 -421 665
rect 1487 631 1583 665
rect -517 569 -483 631
rect -92 563 -26 579
rect -92 529 -76 563
rect -42 529 -26 563
rect -92 513 -26 529
rect 1549 569 1583 631
rect -231 470 -131 486
rect -335 421 -269 437
rect -335 387 -319 421
rect -285 387 -269 421
rect -231 436 -215 470
rect -181 436 -131 470
rect -231 420 -131 436
rect -335 371 -269 387
rect -449 305 -331 321
rect -449 271 -433 305
rect -399 271 -331 305
rect -449 255 -331 271
rect -277 173 -243 337
rect -293 157 -227 173
rect -293 123 -277 157
rect -243 123 -227 157
rect -165 134 -131 420
rect -293 107 -227 123
rect -365 49 -299 65
rect 13 49 47 470
rect -483 0 -407 16
rect -423 -200 -407 0
rect -365 15 -349 49
rect -315 15 47 49
rect 86 49 152 65
rect 86 15 102 49
rect 136 15 152 49
rect -365 -1 -299 15
rect 86 -1 152 15
rect -483 -216 -407 -200
rect -165 -169 -131 -44
rect 13 -60 47 -44
rect 191 -60 225 470
rect 369 335 403 486
rect 369 319 471 335
rect 369 285 421 319
rect 455 285 471 319
rect 369 269 471 285
rect 369 118 403 269
rect 915 66 981 82
rect 264 49 330 65
rect 264 15 280 49
rect 314 15 330 49
rect 915 32 931 66
rect 965 32 981 66
rect 915 16 981 32
rect 1517 60 1549 76
rect 264 -1 330 15
rect 13 -94 191 -60
rect 13 -110 47 -94
rect -92 -169 -26 -153
rect -165 -203 -76 -169
rect -42 -203 -26 -169
rect -92 -219 -26 -203
rect 86 -169 152 -153
rect 86 -203 102 -169
rect 136 -203 152 -169
rect 86 -219 152 -203
rect -517 -742 -483 -680
rect -165 -657 -131 -262
rect 13 -598 47 -262
rect 191 -598 225 -94
rect 280 -153 314 -1
rect 931 -110 965 16
rect 1517 -100 1533 60
rect 1517 -116 1549 -100
rect 264 -169 330 -153
rect 264 -203 280 -169
rect 314 -203 330 -169
rect 264 -219 330 -203
rect 369 -397 403 -246
rect 369 -413 469 -397
rect 369 -447 419 -413
rect 453 -447 469 -413
rect 369 -463 469 -447
rect 573 -413 639 -397
rect 573 -447 589 -413
rect 623 -447 639 -413
rect 573 -463 639 -447
rect 369 -614 403 -463
rect 86 -657 152 -641
rect 489 -657 555 -641
rect -165 -691 102 -657
rect 136 -691 505 -657
rect 539 -691 555 -657
rect 86 -707 152 -691
rect 489 -707 555 -691
rect 1449 -708 1515 -642
rect 1549 -742 1583 -680
rect -517 -776 -421 -742
rect 1487 -776 1583 -742
<< viali >>
rect 178 2473 238 2533
rect 102 2111 136 2145
rect 573 2111 607 2146
rect -476 1510 -416 1570
rect -76 1581 -42 1615
rect 489 1867 523 1901
rect 421 1581 455 1615
rect 191 1471 225 1505
rect -426 1363 -392 1397
rect -349 1247 -315 1281
rect -249 1279 -215 1313
rect -321 986 -287 1020
rect -215 968 -181 1002
rect 102 1363 136 1397
rect 908 1532 942 1566
rect 1086 1532 1120 1566
rect 280 1363 314 1397
rect 997 1389 1031 1423
rect 1563 1360 1579 1560
rect 1579 1360 1597 1560
rect -76 829 -42 863
rect -76 529 -42 563
rect -319 387 -285 421
rect -215 436 -181 470
rect -433 271 -399 305
rect -277 123 -243 157
rect -483 -200 -423 0
rect -349 15 -315 49
rect 102 15 136 49
rect 421 285 455 319
rect 280 15 314 49
rect 931 32 965 66
rect 191 -94 225 -60
rect -76 -203 -42 -169
rect 102 -203 136 -169
rect 1533 -100 1549 60
rect 1549 -100 1567 60
rect 280 -203 314 -169
rect 419 -447 453 -413
rect 589 -447 623 -413
rect 102 -691 136 -657
rect 505 -691 539 -657
rect 842 -692 876 -658
rect 1020 -692 1054 -658
<< metal1 >>
rect 166 2533 250 2539
rect 166 2473 178 2533
rect 238 2473 250 2533
rect 166 2467 250 2473
rect 158 2351 258 2358
rect 158 2348 178 2351
rect 89 2298 178 2348
rect 158 2295 178 2298
rect 238 2295 258 2351
rect 158 2288 258 2295
rect 86 2154 152 2161
rect 567 2155 613 2158
rect 62 2102 72 2154
rect 124 2146 152 2154
rect 554 2146 564 2155
rect 124 2145 564 2146
rect 136 2111 564 2145
rect 124 2102 152 2111
rect 554 2102 564 2111
rect 616 2102 626 2155
rect 86 2095 152 2102
rect 567 2099 613 2102
rect 473 1910 539 1917
rect 473 1858 487 1910
rect 539 1858 549 1910
rect 473 1851 539 1858
rect -92 1615 -26 1631
rect 405 1624 471 1631
rect 405 1615 419 1624
rect -92 1581 -76 1615
rect -42 1581 419 1615
rect -488 1570 -404 1576
rect -488 1510 -476 1570
rect -416 1510 -404 1570
rect -92 1565 -26 1581
rect 405 1572 419 1581
rect 471 1572 481 1624
rect 405 1565 471 1572
rect 892 1566 958 1582
rect 1070 1566 1136 1582
rect 751 1532 908 1566
rect 942 1532 1086 1566
rect 1120 1532 1136 1566
rect 1557 1560 1603 1572
rect -488 1504 -404 1510
rect 175 1514 241 1521
rect 175 1462 182 1514
rect 234 1462 241 1514
rect 175 1455 241 1462
rect 751 1429 785 1532
rect 892 1516 958 1532
rect 1070 1516 1136 1532
rect 981 1432 1047 1439
rect -442 1406 -376 1413
rect 86 1406 152 1413
rect -445 1354 -435 1406
rect -383 1354 -373 1406
rect 62 1354 72 1406
rect 124 1397 152 1406
rect 136 1363 152 1397
rect 124 1354 152 1363
rect -442 1347 -376 1354
rect 86 1347 152 1354
rect 264 1397 330 1413
rect 731 1397 804 1429
rect 264 1363 280 1397
rect 314 1363 804 1397
rect 981 1380 988 1432
rect 1040 1380 1047 1432
rect 981 1373 1047 1380
rect 264 1347 330 1363
rect 1544 1360 1554 1560
rect 1606 1360 1616 1560
rect 1557 1348 1603 1360
rect -365 1290 -299 1297
rect -368 1238 -358 1290
rect -306 1238 -296 1290
rect -268 1270 -258 1322
rect -206 1270 -196 1322
rect -365 1231 -299 1238
rect -337 1020 -271 1036
rect -337 986 -321 1020
rect -287 986 -271 1020
rect -231 1011 -165 1018
rect -337 970 -271 986
rect -234 959 -224 1011
rect -172 959 -162 1011
rect -231 952 -165 959
rect -92 872 -26 879
rect -95 820 -85 872
rect -33 820 -23 872
rect -92 813 -26 820
rect -92 572 -26 579
rect -95 520 -85 572
rect -33 520 -23 572
rect -92 513 -26 520
rect -231 479 -165 486
rect -335 421 -269 437
rect -234 427 -224 479
rect -172 427 -162 479
rect -335 387 -319 421
rect -285 387 -269 421
rect -231 420 -165 427
rect -335 371 -269 387
rect -449 314 -383 321
rect -452 262 -442 314
rect -390 262 -380 314
rect 402 276 412 328
rect 464 276 474 328
rect -449 255 -383 262
rect -293 166 -227 173
rect -296 114 -286 166
rect -234 114 -224 166
rect -293 107 -227 114
rect -365 58 -299 65
rect -489 0 -417 12
rect -368 6 -358 58
rect -306 6 -296 58
rect 86 49 152 65
rect 86 15 102 49
rect 136 15 152 49
rect -493 -200 -483 0
rect -423 -200 -413 0
rect -365 -1 -299 6
rect 86 -1 152 15
rect 264 49 330 65
rect 264 15 280 49
rect 314 15 330 49
rect 912 23 922 75
rect 974 23 984 75
rect 1527 60 1573 72
rect 264 -1 330 15
rect 102 -153 136 -1
rect 175 -51 241 -44
rect 175 -103 182 -51
rect 234 -103 241 -51
rect 175 -110 241 -103
rect 280 -153 314 -1
rect 1523 -100 1533 60
rect 1585 -100 1595 60
rect 1527 -112 1573 -100
rect -92 -160 -26 -153
rect -489 -212 -417 -200
rect -95 -212 -85 -160
rect -33 -212 -23 -160
rect 86 -169 152 -153
rect 86 -203 102 -169
rect 136 -203 152 -169
rect -92 -219 -26 -212
rect 86 -219 152 -203
rect 264 -169 330 -153
rect 1446 -160 1518 -153
rect 1446 -169 1456 -160
rect 264 -203 280 -169
rect 314 -203 1456 -169
rect 264 -219 330 -203
rect 1446 -212 1456 -203
rect 1508 -212 1518 -160
rect 1446 -219 1518 -212
rect 102 -641 136 -219
rect 403 -413 469 -397
rect 573 -404 639 -397
rect 570 -413 580 -404
rect 403 -447 419 -413
rect 453 -447 580 -413
rect 403 -463 469 -447
rect 570 -456 580 -447
rect 632 -456 642 -404
rect 573 -463 639 -456
rect 86 -657 152 -641
rect 489 -648 555 -641
rect 486 -657 496 -648
rect 86 -691 102 -657
rect 136 -691 496 -657
rect 86 -707 152 -691
rect 486 -701 496 -691
rect 548 -701 558 -648
rect 826 -658 892 -642
rect 1004 -658 1070 -642
rect 826 -692 842 -658
rect 876 -692 1020 -658
rect 1054 -692 1499 -658
rect 489 -707 555 -701
rect 826 -708 892 -692
rect 1004 -708 1070 -692
<< via1 >>
rect 178 2473 238 2533
rect 178 2295 238 2351
rect 72 2145 124 2154
rect 564 2146 616 2155
rect 72 2111 102 2145
rect 102 2111 124 2145
rect 564 2111 573 2146
rect 573 2111 607 2146
rect 607 2111 616 2146
rect 72 2102 124 2111
rect 564 2102 616 2111
rect 487 1901 539 1910
rect 487 1867 489 1901
rect 489 1867 523 1901
rect 523 1867 539 1901
rect 487 1858 539 1867
rect 419 1615 471 1624
rect 419 1581 421 1615
rect 421 1581 455 1615
rect 455 1581 471 1615
rect -476 1510 -416 1570
rect 419 1572 471 1581
rect 182 1505 234 1514
rect 182 1471 191 1505
rect 191 1471 225 1505
rect 225 1471 234 1505
rect 182 1462 234 1471
rect -435 1397 -383 1406
rect -435 1363 -426 1397
rect -426 1363 -392 1397
rect -392 1363 -383 1397
rect -435 1354 -383 1363
rect 72 1397 124 1406
rect 72 1363 102 1397
rect 102 1363 124 1397
rect 72 1354 124 1363
rect 988 1423 1040 1432
rect 988 1389 997 1423
rect 997 1389 1031 1423
rect 1031 1389 1040 1423
rect 988 1380 1040 1389
rect 1554 1360 1563 1560
rect 1563 1360 1597 1560
rect 1597 1360 1606 1560
rect -358 1281 -306 1290
rect -358 1247 -349 1281
rect -349 1247 -315 1281
rect -315 1247 -306 1281
rect -358 1238 -306 1247
rect -258 1313 -206 1322
rect -258 1279 -249 1313
rect -249 1279 -215 1313
rect -215 1279 -206 1313
rect -258 1270 -206 1279
rect -224 1002 -172 1011
rect -224 968 -215 1002
rect -215 968 -181 1002
rect -181 968 -172 1002
rect -224 959 -172 968
rect -85 863 -33 872
rect -85 829 -76 863
rect -76 829 -42 863
rect -42 829 -33 863
rect -85 820 -33 829
rect -85 563 -33 572
rect -85 529 -76 563
rect -76 529 -42 563
rect -42 529 -33 563
rect -85 520 -33 529
rect -224 470 -172 479
rect -224 436 -215 470
rect -215 436 -181 470
rect -181 436 -172 470
rect -224 427 -172 436
rect -442 305 -390 314
rect -442 271 -433 305
rect -433 271 -399 305
rect -399 271 -390 305
rect -442 262 -390 271
rect 412 319 464 328
rect 412 285 421 319
rect 421 285 455 319
rect 455 285 464 319
rect 412 276 464 285
rect -286 157 -234 166
rect -286 123 -277 157
rect -277 123 -243 157
rect -243 123 -234 157
rect -286 114 -234 123
rect -358 49 -306 58
rect -358 15 -349 49
rect -349 15 -315 49
rect -315 15 -306 49
rect -358 6 -306 15
rect -483 -200 -423 0
rect 922 66 974 75
rect 922 32 931 66
rect 931 32 965 66
rect 965 32 974 66
rect 922 23 974 32
rect 182 -60 234 -51
rect 182 -94 191 -60
rect 191 -94 225 -60
rect 225 -94 234 -60
rect 182 -103 234 -94
rect 1533 -100 1567 60
rect 1567 -100 1585 60
rect -85 -169 -33 -160
rect -85 -203 -76 -169
rect -76 -203 -42 -169
rect -42 -203 -33 -169
rect -85 -212 -33 -203
rect 1456 -212 1508 -160
rect 580 -413 632 -404
rect 580 -447 589 -413
rect 589 -447 623 -413
rect 623 -447 632 -413
rect 580 -456 632 -447
rect 496 -657 548 -648
rect 496 -691 505 -657
rect 505 -691 539 -657
rect 539 -691 548 -657
rect 496 -701 548 -691
<< metal2 >>
rect 158 2533 258 2543
rect 158 2473 178 2533
rect 238 2473 258 2533
rect 158 2351 258 2473
rect 158 2295 178 2351
rect 238 2295 258 2351
rect 72 2154 124 2164
rect -476 1570 -416 1580
rect -476 1500 -416 1510
rect -435 1406 -383 1416
rect -435 1344 -383 1354
rect 72 1406 124 2102
rect 158 1516 258 2295
rect 564 2155 616 2165
rect 564 2092 616 2102
rect 487 1910 539 1920
rect 487 1848 539 1858
rect 419 1624 471 1634
rect 419 1562 471 1572
rect 158 1460 180 1516
rect 236 1460 258 1516
rect 158 1438 258 1460
rect 72 1344 124 1354
rect -426 324 -392 1344
rect -260 1324 -204 1334
rect -358 1290 -306 1300
rect -260 1258 -204 1268
rect -358 1228 -306 1238
rect -442 314 -390 324
rect -442 252 -390 262
rect -358 68 -324 1228
rect -224 1011 -172 1021
rect -224 949 -172 959
rect -215 489 -181 949
rect -85 872 -33 882
rect -85 810 -33 820
rect -76 582 -42 810
rect -85 572 -33 582
rect -85 510 -33 520
rect -224 479 -172 489
rect -224 417 -172 427
rect -288 168 -232 178
rect -288 102 -232 112
rect -358 58 -306 68
rect -483 0 -423 10
rect -358 -4 -306 6
rect -76 -150 -42 510
rect 437 338 471 1562
rect 412 328 471 338
rect 464 276 471 328
rect 412 266 471 276
rect 171 -49 245 -40
rect 171 -105 180 -49
rect 236 -105 245 -49
rect 171 -114 245 -105
rect -483 -210 -423 -200
rect -85 -160 -33 -150
rect -85 -222 -33 -212
rect 505 -638 539 1848
rect 573 -394 607 2092
rect 1552 1560 1608 1570
rect 977 1434 1051 1439
rect 977 1378 986 1434
rect 1042 1378 1051 1434
rect 977 1373 1051 1378
rect 1552 1350 1608 1360
rect 920 77 976 87
rect 920 11 976 21
rect 1533 60 1589 70
rect 1533 -110 1589 -100
rect 1456 -160 1508 -150
rect 1456 -222 1508 -212
rect 573 -404 632 -394
rect 573 -456 580 -404
rect 573 -466 632 -456
rect 496 -648 548 -638
rect 496 -711 548 -701
<< via2 >>
rect -476 1510 -416 1570
rect 180 1514 236 1516
rect 180 1462 182 1514
rect 182 1462 234 1514
rect 234 1462 236 1514
rect 180 1460 236 1462
rect -260 1322 -204 1324
rect -260 1270 -258 1322
rect -258 1270 -206 1322
rect -206 1270 -204 1322
rect -260 1268 -204 1270
rect -288 166 -232 168
rect -288 114 -286 166
rect -286 114 -234 166
rect -234 114 -232 166
rect -288 112 -232 114
rect -483 -200 -423 0
rect 180 -51 236 -49
rect 180 -103 182 -51
rect 182 -103 234 -51
rect 234 -103 236 -51
rect 180 -105 236 -103
rect 986 1432 1042 1434
rect 986 1380 988 1432
rect 988 1380 1040 1432
rect 1040 1380 1042 1432
rect 986 1378 1042 1380
rect 1552 1360 1554 1560
rect 1554 1360 1606 1560
rect 1606 1360 1608 1560
rect 920 75 976 77
rect 920 23 922 75
rect 922 23 974 75
rect 974 23 976 75
rect 920 21 976 23
rect 1533 -100 1585 60
rect 1585 -100 1589 60
<< metal3 >>
rect -1000 1570 2140 1700
rect -1000 1510 -476 1570
rect -416 1560 2140 1570
rect -416 1516 1552 1560
rect -416 1510 180 1516
rect -1000 1460 180 1510
rect 236 1460 1552 1516
rect -1000 1434 1552 1460
rect -1000 1378 986 1434
rect 1042 1378 1552 1434
rect -1000 1360 1552 1378
rect 1608 1360 2140 1560
rect -1000 1324 2140 1360
rect -1000 1300 -260 1324
rect -270 1268 -260 1300
rect -204 1300 2140 1324
rect -204 1268 -194 1300
rect -270 1263 -194 1268
rect -298 168 -222 173
rect -298 112 -288 168
rect -232 112 -222 168
rect -298 100 -222 112
rect -1000 77 2140 100
rect -1000 21 920 77
rect 976 60 2140 77
rect 976 21 1533 60
rect -1000 0 1533 21
rect -1000 -200 -483 0
rect -423 -49 1533 0
rect -423 -105 180 -49
rect 236 -100 1533 -49
rect 1589 -100 2140 60
rect 236 -105 2140 -100
rect -423 -200 2140 -105
rect -1000 -300 2140 -200
use bias2  x2
timestamp 1731242581
transform 1 0 939 0 1 633
box -902 -1344 608 1777
use sky130_fd_pr__nfet_01v8_ZJWC73  XM1
timestamp 1729864714
transform 1 0 119 0 -1 302
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_ZJWC73  XM2
timestamp 1729864714
transform 1 0 -59 0 -1 302
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_ZJWC73  XM3
timestamp 1729864714
transform 1 0 -59 0 -1 -430
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_ZJWC73  XM4
timestamp 1729864714
transform 1 0 119 0 -1 -430
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_PU4Y8N  XM5
timestamp 1729864714
transform 1 0 -304 0 1 288
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_AH2TBC  XM6
timestamp 1729864714
transform 1 0 119 0 1 1136
box -154 -242 154 242
use sky130_fd_pr__pfet_01v8_AH2TBC  XM7
timestamp 1729864714
transform 1 0 -59 0 1 1868
box -154 -242 154 242
use sky130_fd_pr__pfet_01v8_AH2TBC  XM8
timestamp 1729864714
transform 1 0 -59 0 1 1136
box -154 -242 154 242
use sky130_fd_pr__pfet_01v8_AH2TBC  XM9
timestamp 1729864714
transform 1 0 119 0 1 1868
box -154 -242 154 242
use sky130_fd_pr__pfet_01v8_58PGBE  XM10
timestamp 1729864714
transform 1 0 -304 0 1 1136
box -109 -122 109 122
use sky130_fd_pr__nfet_01v8_4NLQMD  XM11
timestamp 1729864714
transform 1 0 -59 0 1 -77
box -118 -71 118 71
use sky130_fd_pr__pfet_01v8_W2SF2B  XM12
timestamp 1729864714
transform 1 0 -59 0 1 1489
box -154 -107 154 107
use sky130_fd_pr__pfet_01v8_AH2TBC  XM13
timestamp 1729864714
transform -1 0 297 0 1 1136
box -154 -242 154 242
use sky130_fd_pr__nfet_01v8_ZJWC73  XM14
timestamp 1729864714
transform -1 0 297 0 1 302
box -118 -206 118 206
use sky130_fd_pr__nfet_01v8_ZJWC73  XM15
timestamp 1729864714
transform -1 0 297 0 1 -430
box -118 -206 118 206
use sky130_fd_pr__pfet_01v8_AH2TBC  XM16
timestamp 1729864714
transform -1 0 297 0 1 1868
box -154 -242 154 242
<< labels >>
flabel metal3 -1000 1482 -966 1518 0 FreeSans 320 0 0 0 vdd
flabel metal3 -1000 -118 -966 -82 0 FreeSans 320 0 0 0 vss
port 1 nsew
flabel metal1 -319 387 -285 421 0 FreeSans 320 0 0 0 upb
port 2 nsew
flabel metal1 -321 986 -287 1020 0 FreeSans 320 0 0 0 down
port 3 nsew
flabel metal2 -215 702 -181 736 0 FreeSans 320 0 0 0 out
port 4 nsew
<< end >>
