magic
tech sky130A
magscale 1 2
timestamp 1726263301
<< nwell >>
rect 6 991 40 1005
rect 198 991 232 1005
rect -40 961 278 991
rect 6 953 40 961
rect 198 953 232 961
rect 294 953 328 999
rect -90 811 -56 845
rect 102 811 136 845
rect 294 811 328 845
rect 376 669 630 850
<< pwell >>
rect 696 426 3735 453
rect -170 298 3735 426
rect 61 212 147 298
<< poly >>
rect -106 1190 -40 1206
rect -106 1156 -90 1190
rect -56 1188 -40 1190
rect 86 1190 152 1206
rect -56 1173 -10 1188
rect 86 1173 102 1190
rect -56 1156 102 1173
rect 136 1173 152 1190
rect 278 1190 344 1206
rect 278 1173 294 1190
rect 136 1156 294 1173
rect 328 1156 344 1190
rect -106 1143 344 1156
rect -106 1140 -10 1143
rect -40 994 -10 1140
rect 56 1140 182 1143
rect 56 994 86 1140
rect 152 994 182 1140
rect 248 1140 344 1143
rect 248 994 278 1140
rect -40 964 278 994
rect -40 898 -10 964
rect 56 898 86 964
rect 152 898 182 964
rect 248 898 278 964
rect 42 530 126 540
rect -86 500 -20 516
rect -86 466 -70 500
rect -36 466 -20 500
rect 42 496 58 530
rect 92 496 126 530
rect 42 484 126 496
rect 42 480 606 484
rect -86 412 -20 466
rect 76 438 606 480
rect 96 412 126 438
<< polycont >>
rect -90 1156 -56 1190
rect 102 1156 136 1190
rect 294 1156 328 1190
rect -70 466 -36 500
rect 58 496 92 530
<< locali >>
rect 6 1620 62 1638
rect 6 1586 22 1620
rect 56 1586 62 1620
rect 6 1568 62 1586
rect 198 1621 232 1639
rect 198 1587 206 1621
rect 198 1586 516 1587
rect -106 1190 -40 1206
rect -106 1156 -90 1190
rect -56 1156 -40 1190
rect -106 1140 -40 1156
rect -90 1097 -56 1140
rect -158 1005 -56 1097
rect -158 416 -124 1005
rect -90 811 -56 900
rect 6 897 40 1568
rect 86 1190 152 1206
rect 86 1156 102 1190
rect 136 1156 152 1190
rect 86 1140 152 1156
rect 102 1113 136 1140
rect 102 811 136 900
rect 198 897 232 1586
rect 278 1190 344 1206
rect 278 1156 294 1190
rect 328 1156 344 1190
rect 278 1140 344 1156
rect 294 1113 328 1140
rect 1402 959 1926 974
rect 1402 925 1585 959
rect 1619 925 1677 959
rect 1711 925 1769 959
rect 1803 925 1861 959
rect 1895 925 1926 959
rect 294 811 328 900
rect 1402 811 1926 925
rect -90 777 -40 811
rect -6 777 52 811
rect 86 777 144 811
rect 178 777 236 811
rect 270 777 651 811
rect 3629 777 3646 811
rect 42 530 108 540
rect -86 500 -20 516
rect -86 466 -70 500
rect -36 466 -20 500
rect 42 496 58 530
rect 92 496 108 530
rect 3252 514 3352 530
rect 42 480 108 496
rect 142 480 542 511
rect 576 480 718 511
rect -86 450 -20 466
rect 142 464 718 480
rect 966 464 1099 511
rect 1347 464 1480 511
rect 1728 464 1861 511
rect 2109 464 2242 511
rect 2490 464 2623 511
rect 2871 464 3004 511
rect 3252 480 3302 514
rect 3336 513 3352 514
rect 3563 514 3629 530
rect 3336 480 3460 513
rect 3563 505 3579 514
rect 3252 465 3460 480
rect 3517 480 3579 505
rect 3613 480 3629 514
rect 3517 471 3629 480
rect 3252 464 3352 465
rect 3563 464 3629 471
rect -158 308 -98 416
rect 46 267 80 363
rect 142 361 176 464
rect 334 416 368 464
rect 526 416 560 464
rect 238 267 272 367
rect 430 267 464 367
rect 622 267 656 367
rect 46 233 87 267
rect 121 233 179 267
rect 213 233 271 267
rect 305 233 363 267
rect 397 233 455 267
rect 489 233 547 267
rect 581 233 639 267
rect 3318 233 3353 267
rect 3629 233 3646 267
<< viali >>
rect 22 1586 56 1620
rect 206 1587 240 1621
rect 298 1587 332 1621
rect 390 1587 424 1621
rect 482 1587 516 1621
rect 1585 925 1619 959
rect 1677 925 1711 959
rect 1769 925 1803 959
rect 1861 925 1895 959
rect -40 777 -6 811
rect 52 777 86 811
rect 144 777 178 811
rect 236 777 270 811
rect -70 466 -36 500
rect 58 496 92 530
rect 542 480 576 514
rect 3302 480 3336 514
rect 3579 480 3613 514
rect 87 233 121 267
rect 179 233 213 267
rect 271 233 305 267
rect 363 233 397 267
rect 455 233 489 267
rect 547 233 581 267
rect 639 233 673 267
<< metal1 >>
rect 3353 1651 3629 1652
rect -158 1621 3629 1651
rect -158 1620 206 1621
rect -158 1586 22 1620
rect 56 1587 206 1620
rect 240 1587 298 1621
rect 332 1587 390 1621
rect 424 1587 482 1621
rect 516 1587 3629 1621
rect 56 1586 3629 1587
rect -158 1555 3629 1586
rect 414 1181 506 1555
rect 1402 959 1926 974
rect 1402 925 1585 959
rect 1619 925 1677 959
rect 1711 925 1769 959
rect 1803 925 1861 959
rect 1895 925 1926 959
rect 1402 842 1926 925
rect 3353 842 3629 1555
rect -90 811 3318 842
rect -90 777 -40 811
rect -6 777 52 811
rect 86 777 144 811
rect 178 777 236 811
rect 270 777 3318 811
rect -90 746 3318 777
rect 3629 746 3646 842
rect -158 564 108 630
rect 42 530 108 564
rect -158 500 -20 516
rect -158 466 -70 500
rect -36 466 -20 500
rect 42 496 58 530
rect 92 496 108 530
rect 42 480 108 496
rect 526 514 3352 530
rect 526 480 542 514
rect 576 480 3302 514
rect 3336 480 3352 514
rect -158 450 -20 466
rect 526 464 3352 480
rect 3563 514 3629 530
rect 3563 480 3579 514
rect 3613 480 3629 514
rect 3563 464 3629 480
rect -158 297 3353 298
rect -158 267 3417 297
rect -158 233 87 267
rect 121 233 179 267
rect 213 233 271 267
rect 305 233 363 267
rect 397 233 455 267
rect 489 233 547 267
rect 581 233 639 267
rect 673 233 3417 267
rect -158 202 3417 233
rect 3629 202 3646 298
use tap_1_gnd  sky130_fd_sc_hd__tapvgnd_1_0
timestamp 1726262061
transform 1 0 58 0 -1 250
box 0 -48 92 195
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 3646 0 1 250
box -38 -48 130 592
use tap_1_pwr  tap_1_pwr_0
timestamp 1726200578
transform 1 0 414 0 1 589
box -38 261 130 592
use inv_0p25  x1
timestamp 1726261667
transform -1 0 1121 0 -1 12
box -313 -837 110 -190
use inv_0p25  x2
timestamp 1726261667
transform -1 0 1502 0 -1 12
box -313 -837 110 -190
use inv_0p25  x3
timestamp 1726261667
transform -1 0 1883 0 -1 12
box -313 -837 110 -190
use inv_0p25  x4
timestamp 1726261667
transform -1 0 2264 0 -1 12
box -313 -837 110 -190
use inv_0p25  x5
timestamp 1726261667
transform -1 0 2645 0 -1 12
box -313 -837 110 -190
use sky130_fd_sc_hd__inv_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715908107
transform 1 0 3353 0 1 250
box -38 -48 314 592
use inv_0p25  x12
timestamp 1726261667
transform -1 0 740 0 -1 12
box -313 -837 110 -190
use inv_0p25  x13
timestamp 1726261667
transform -1 0 3026 0 -1 12
box -313 -837 110 -190
use sky130_fd_pr__nfet_01v8_NAAUVB  XM1
timestamp 1726197802
transform 1 0 -26 0 1 362
box -118 -76 118 76
use sky130_fd_pr__pfet_01v8_52X2FE  XM2
timestamp 1726197802
transform 1 0 119 0 -1 1059
box -257 -112 257 112
use sky130_fd_pr__pfet_01v8_52X2FE  XM3
timestamp 1726197802
transform 1 0 119 0 -1 899
box -257 -112 257 112
use sky130_fd_pr__nfet_01v8_YEG85W  XM4
timestamp 1726197802
transform 1 0 351 0 1 362
box -317 -76 317 76
use sky130_fd_pr__res_xhigh_po_0p35_JAND4E  XR3
timestamp 1726197802
transform 0 1 1040 -1 0 1272
box -367 -886 367 886
<< labels >>
flabel metal1 -158 1555 -62 1651 0 FreeSans 320 0 0 0 vdd
port 0 nsew
flabel metal1 3533 1556 3629 1652 0 FreeSans 320 0 0 0 vdd
port 1 nsew
flabel metal1 -158 202 -62 298 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal1 -158 450 -92 516 0 FreeSans 240 0 0 0 vctrl
port 5 nsew
flabel metal1 -158 564 -92 630 0 FreeSans 240 0 0 0 vstart
port 6 nsew
flabel metal1 3563 464 3629 530 0 FreeSans 240 0 0 0 vo
port 7 nsew
flabel metal1 3533 202 3629 297 0 FreeSans 320 0 0 0 vss
port 3 nsew
<< end >>
