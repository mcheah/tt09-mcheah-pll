magic
tech sky130A
magscale 1 2
timestamp 1731242581
<< pwell >>
rect 2319 4826 2405 4923
<< metal1 >>
rect 2310 4911 2414 4933
rect 2310 4859 2336 4911
rect 2388 4859 2414 4911
rect 2310 4837 2414 4859
rect -229 4758 280 4764
rect -229 4652 -219 4758
rect 268 4652 280 4758
rect -229 4646 280 4652
rect 4328 4758 4905 4764
rect 4328 4652 4340 4758
rect 4895 4652 4905 4758
rect 4328 4646 4905 4652
<< via1 >>
rect 2336 4859 2388 4911
rect -219 4652 268 4758
rect 4340 4652 4895 4758
<< metal2 >>
rect 2310 4913 2414 4933
rect 2310 4857 2334 4913
rect 2390 4857 2414 4913
rect 2310 4837 2414 4857
rect -236 4758 285 4774
rect -236 4652 -220 4758
rect 268 4652 285 4758
rect -236 4636 285 4652
rect 4323 4758 4912 4774
rect 4323 4652 4340 4758
rect 4896 4652 4912 4758
rect 4323 4636 4912 4652
<< via2 >>
rect 2334 4911 2390 4913
rect 2334 4859 2336 4911
rect 2336 4859 2388 4911
rect 2388 4859 2390 4911
rect 2334 4857 2390 4859
rect -220 4652 -219 4758
rect -219 4652 -156 4758
rect 4824 4652 4895 4758
rect 4895 4652 4896 4758
<< metal3 >>
rect 2310 4917 2414 4933
rect 2310 4853 2330 4917
rect 2394 4853 2414 4917
rect 2310 4837 2414 4853
rect -236 4758 -140 4774
rect -236 4652 -220 4758
rect -156 4652 -140 4758
rect -236 4504 -140 4652
rect 4808 4758 4912 4774
rect 4808 4652 4824 4758
rect 4896 4652 4912 4758
rect 4808 4516 4912 4652
rect 4808 -240 4920 0
rect 4800 -9484 4920 -240
<< via3 >>
rect 2330 4913 2394 4917
rect 2330 4857 2334 4913
rect 2334 4857 2390 4913
rect 2390 4857 2394 4913
rect 2330 4853 2394 4857
<< metal4 >>
rect 2310 4917 2414 4933
rect 2310 4853 2330 4917
rect 2394 4853 2414 4917
rect 2310 4437 2414 4853
rect 2310 -9856 2414 183
use tap_1_gnd  tap_1_gnd_0
timestamp 1726262061
transform 1 0 2316 0 1 4885
box 0 -48 92 195
use sky130_fd_pr__cap_mim_m3_1_P73DWX  XC1
timestamp 1731188831
transform -1 0 2164 0 1 2258
box -2404 -2258 2404 2258
use sky130_fd_pr__cap_mim_m3_1_PX3DWX  XC2
timestamp 1731188749
transform 1 0 7212 0 1 -7254
box -7108 -2602 2404 11890
use sky130_fd_pr__res_high_po_0p69_T6VK6H  XR1
timestamp 1730848472
transform 0 1 2304 -1 0 4705
box -121 -2503 121 2503
<< labels >>
flabel metal4 2310 -9856 2406 -9760 0 FreeSans 320 0 0 0 vss
port 1 nsew
flabel metal3 -236 4657 -140 4753 0 FreeSans 320 0 0 0 in
port 0 nsew
<< end >>
