magic
tech sky130A
magscale 1 2
timestamp 1731188749
<< metal3 >>
rect -2404 11770 -2300 11890
rect -2404 11742 2404 11770
rect -2404 7282 -2384 11742
rect -2320 7282 2404 11742
rect -2404 7254 2404 7282
rect -7108 6986 2404 7014
rect -7108 2526 -2384 6986
rect -2320 2526 2404 6986
rect -7108 2498 2404 2526
rect -7108 2230 2404 2258
rect -7108 -2230 -2384 2230
rect -2320 -2230 2404 2230
rect -7108 -2258 2404 -2230
<< via3 >>
rect -2384 7282 -2320 11742
rect -2384 2526 -2320 6986
rect -2384 -2230 -2320 2230
<< mimcap >>
rect -2072 11690 2364 11730
rect -2072 7334 -2032 11690
rect 2324 7334 2364 11690
rect -2072 7294 2364 7334
rect -7068 6934 -2632 6974
rect -7068 2578 -7028 6934
rect -2672 2578 -2632 6934
rect -7068 2538 -2632 2578
rect -2072 6934 2364 6974
rect -2072 2578 -2032 6934
rect 2324 2578 2364 6934
rect -2072 2538 2364 2578
rect -7068 2178 -2632 2218
rect -7068 -2178 -7028 2178
rect -2672 -2178 -2632 2178
rect -7068 -2218 -2632 -2178
rect -2072 2178 2364 2218
rect -2072 -2178 -2032 2178
rect 2324 -2178 2364 2178
rect -2072 -2218 2364 -2178
<< mimcapcontact >>
rect -2032 7334 2324 11690
rect -7028 2578 -2672 6934
rect -2032 2578 2324 6934
rect -7028 -2178 -2672 2178
rect -2032 -2178 2324 2178
<< metal4 >>
rect -2404 11742 -2300 11770
rect -4902 6935 -4798 7334
rect -2404 7282 -2384 11742
rect -2320 7282 -2300 11742
rect 94 11691 198 11890
rect -2033 11690 2325 11691
rect -2033 7334 -2032 11690
rect 2324 7334 2325 11690
rect -2033 7333 2325 7334
rect -2404 6986 -2300 7282
rect -7029 6934 -2671 6935
rect -7029 2578 -7028 6934
rect -2672 2578 -2671 6934
rect -7029 2577 -2671 2578
rect -4902 2179 -4798 2577
rect -2404 2526 -2384 6986
rect -2320 2526 -2300 6986
rect 94 6935 198 7333
rect -2033 6934 2325 6935
rect -2033 2578 -2032 6934
rect 2324 2578 2325 6934
rect -2033 2577 2325 2578
rect -2404 2230 -2300 2526
rect -7029 2178 -2671 2179
rect -7029 -2178 -7028 2178
rect -2672 -2178 -2671 2178
rect -7029 -2179 -2671 -2178
rect -4902 -2498 -4798 -2179
rect -2404 -2230 -2384 2230
rect -2320 -2230 -2300 2230
rect 94 2179 198 2577
rect -2033 2178 2325 2179
rect -2033 -2178 -2032 2178
rect 2324 -2178 2325 2178
rect -2033 -2179 2325 -2178
rect -2404 -2258 -2300 -2230
rect 94 -2498 198 -2179
rect -4902 -2602 198 -2498
<< labels >>
flabel metal4 -4902 -2602 -4798 -2498 0 FreeSans 320 0 0 0 c1
port 0 nsew
flabel metal3 -2404 11787 -2300 11890 0 FreeSans 320 0 0 0 c0
port 1 nsew
<< properties >>
string FIXED_BBOX -2404 7254 2112 11770
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22.175 l 22.175 val 1.0k carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
